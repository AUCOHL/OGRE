VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
  DATABASE MICRONS 2000 ;
END UNITS

PROPERTYDEFINITIONS
    LAYER LEF58_CORNERSPACING STRING ;
END PROPERTYDEFINITIONS

CLEARANCEMEASURE EUCLIDEAN ;
MANUFACTURINGGRID 0.0005 ;
USEMINSPACING OBS ON ;

LAYER Metal1
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.10 0.10 ;
  WIDTH 0.05 ;
  AREA 0.0115 ;
  MINWIDTH 0.05 ;
  SPACINGTABLE
    PARALLELRUNLENGTH  0.0 0.22 0.47 0.63 1.50
    WIDTH 0.0         0.05 0.05 0.05 0.05 0.05
    WIDTH 0.10        0.05 0.06 0.06 0.06 0.06
    WIDTH 0.28        0.05 0.10 0.10 0.10 0.10
    WIDTH 0.47        0.05 0.10 0.13 0.13 0.13
    WIDTH 0.63        0.05 0.10 0.13 0.15 0.15
    WIDTH 1.50        0.05 0.10 0.13 0.15 0.50 ;
  SPACING 0.06 ENDOFLINE 0.06 WITHIN 0.025 ;
END Metal1

LAYER Via1
  TYPE CUT ;
  SPACING 0.075 ;
  WIDTH 0.05 ;
END Via1

LAYER Metal2
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.10 0.10 ;
  WIDTH 0.05 ;
  AREA 0.014 ;
  MINWIDTH 0.05 ;
  SPACINGTABLE
    PARALLELRUNLENGTH  0.0 0.22 0.47 0.63 1.5
    WIDTH 0.0         0.05 0.05 0.05 0.05 0.05
    WIDTH 0.09        0.05 0.06 0.06 0.06 0.06
    WIDTH 0.16        0.05 0.10 0.10 0.10 0.10
    WIDTH 0.47        0.05 0.10 0.13 0.13 0.13
    WIDTH 0.63        0.05 0.10 0.13 0.15 0.15
    WIDTH 1.5         0.05 0.10 0.13 0.15 0.50 ;
  SPACING 0.08 ENDOFLINE 0.08 WITHIN 0.025 ;
  SPACING 0.10 ENDOFLINE 0.08 WITHIN 0.025 PARALLELEDGE 0.10 WITHIN 0.025 ;
  PROPERTY LEF58_CORNERSPACING "CORNERSPACING CONVEXCORNER EXCEPTEOL 0.08
    WIDTH 0.00 SPACING 0.10
    WIDTH 0.20 SPACING 0.20
    WIDTH 0.50 SPACING 0.30 ;" ;
END Metal2

LAYER Via2
  TYPE CUT ;
  SPACING 0.075 ;
  WIDTH 0.05 ;
  SPACING 0.155 ADJACENTCUTS 3 WITHIN 0.200 ;
END Via2

LAYER Metal3
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.10 0.10 ;
  WIDTH 0.05 ;
  AREA 0.017 ;
  MINWIDTH 0.05 ;
  SPACINGTABLE
    PARALLELRUNLENGTH  0.0 0.22 0.47 0.63 1.5
    WIDTH 0.0         0.05 0.05 0.05 0.05 0.05
    WIDTH 0.09        0.05 0.06 0.06 0.06 0.06
    WIDTH 0.16        0.05 0.10 0.10 0.10 0.10
    WIDTH 0.47        0.05 0.10 0.13 0.13 0.13
    WIDTH 0.63        0.05 0.10 0.13 0.15 0.15
    WIDTH 1.5         0.05 0.10 0.13 0.15 0.50 ;
  SPACING 0.08 ENDOFLINE 0.08 WITHIN 0.025 ;
  SPACING 0.10 ENDOFLINE 0.08 WITHIN 0.025 PARALLELEDGE 0.10 WITHIN 0.025 ;
  PROPERTY LEF58_CORNERSPACING "CORNERSPACING CONVEXCORNER EXCEPTEOL 0.08
    WIDTH 0.00 SPACING 0.10
    WIDTH 0.20 SPACING 0.20
    WIDTH 0.50 SPACING 0.30 ;" ;
END Metal3

LAYER Via3
  TYPE CUT ;
  SPACING 0.075 ;
  WIDTH 0.05 ;
  SPACING 0.155 ADJACENTCUTS 3 WITHIN 0.200 ;
END Via3

LAYER Metal4
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.10 0.10 ;
  WIDTH 0.05 ;
  AREA 0.017 ;
  MINWIDTH 0.05 ;
  SPACINGTABLE
    PARALLELRUNLENGTH  0.0 0.22 0.47 0.63 1.5
    WIDTH 0.0         0.05 0.05 0.05 0.05 0.05
    WIDTH 0.09        0.05 0.06 0.06 0.06 0.06
    WIDTH 0.16        0.05 0.10 0.10 0.10 0.10
    WIDTH 0.47        0.05 0.10 0.13 0.13 0.13
    WIDTH 0.63        0.05 0.10 0.13 0.15 0.15
    WIDTH 1.5         0.05 0.10 0.13 0.15 0.50 ;
  SPACING 0.08 ENDOFLINE 0.08 WITHIN 0.025 ;
  SPACING 0.10 ENDOFLINE 0.08 WITHIN 0.025 PARALLELEDGE 0.10 WITHIN 0.025 ;
  PROPERTY LEF58_CORNERSPACING "CORNERSPACING CONVEXCORNER EXCEPTEOL 0.08
    WIDTH 0.00 SPACING 0.10
    WIDTH 0.20 SPACING 0.20
    WIDTH 0.50 SPACING 0.30 ;" ;
END Metal4

LAYER Via4
  TYPE CUT ;
  SPACING 0.075 ;
  WIDTH 0.05 ;
  SPACING 0.155 ADJACENTCUTS 3 WITHIN 0.200 ;
END Via4

LAYER Metal5
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.10 0.10 ;
  WIDTH 0.05 ;
  AREA 0.017 ;
  MINWIDTH 0.05 ;
  SPACINGTABLE
    PARALLELRUNLENGTH  0.0 0.22 0.47 0.63 1.5
    WIDTH 0.0         0.05 0.05 0.05 0.05 0.05
    WIDTH 0.09        0.05 0.06 0.06 0.06 0.06
    WIDTH 0.16        0.05 0.10 0.10 0.10 0.10
    WIDTH 0.47        0.05 0.10 0.13 0.13 0.13
    WIDTH 0.63        0.05 0.10 0.13 0.15 0.15
    WIDTH 1.5         0.05 0.10 0.13 0.15 0.50 ;
  SPACING 0.08 ENDOFLINE 0.08 WITHIN 0.025 ;
  SPACING 0.10 ENDOFLINE 0.08 WITHIN 0.025 PARALLELEDGE 0.10 WITHIN 0.025 ;
  PROPERTY LEF58_CORNERSPACING "CORNERSPACING CONVEXCORNER EXCEPTEOL 0.08
    WIDTH 0.00 SPACING 0.10
    WIDTH 0.20 SPACING 0.20
    WIDTH 0.50 SPACING 0.30 ;" ;
END Metal5

LAYER Via5
  TYPE CUT ;
  SPACING 0.075 ;
  WIDTH 0.05 ;
  SPACING 0.155 ADJACENTCUTS 3 WITHIN 0.200 ;
END Via5

LAYER Metal6
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.15 0.15 ;
  WIDTH 0.07 ;
  AREA 0.025 ;
  MINWIDTH 0.07 ;
  SPACINGTABLE
    PARALLELRUNLENGTH  0.0 0.22 0.47 0.63 1.5
    WIDTH 0.0         0.08 0.08 0.08 0.08 0.08
    WIDTH 0.10        0.08 0.12 0.12 0.12 0.12
    WIDTH 0.16        0.08 0.12 0.15 0.15 0.15
    WIDTH 0.47        0.08 0.12 0.15 0.18 0.18
    WIDTH 0.63        0.08 0.12 0.15 0.18 0.25
    WIDTH 1.5         0.08 0.12 0.15 0.18 0.50 ;
  SPACING 0.10 ENDOFLINE 0.10 WITHIN 0.035 ;
  SPACING 0.12 ENDOFLINE 0.10 WITHIN 0.035 PARALLELEDGE 0.12 WITHIN 0.035 ;
  PROPERTY LEF58_CORNERSPACING "CORNERSPACING CONVEXCORNER EXCEPTEOL 0.08
    WIDTH 0.00 SPACING 0.10
    WIDTH 0.20 SPACING 0.20
    WIDTH 0.50 SPACING 0.30 ;" ;
END Metal6

LAYER Via6
  TYPE CUT ;
  SPACING 0.10 ;
  WIDTH 0.07 ;
  SPACING 0.20 ADJACENTCUTS 3 WITHIN 0.25 ;
END Via6

LAYER Metal7
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.15 0.15 ;
  WIDTH 0.07 ;
  AREA 0.025 ;
  MINWIDTH 0.07 ;
  SPACINGTABLE
    PARALLELRUNLENGTH  0.0 0.22 0.47 0.63 1.5
    WIDTH 0.0         0.08 0.08 0.08 0.08 0.08
    WIDTH 0.10        0.08 0.12 0.12 0.12 0.12
    WIDTH 0.16        0.08 0.12 0.15 0.15 0.15
    WIDTH 0.47        0.08 0.12 0.15 0.18 0.18
    WIDTH 0.63        0.08 0.12 0.15 0.18 0.25
    WIDTH 1.5         0.08 0.12 0.15 0.18 0.50 ;
  SPACING 0.10 ENDOFLINE 0.10 WITHIN 0.035 ;
  SPACING 0.12 ENDOFLINE 0.10 WITHIN 0.035 PARALLELEDGE 0.12 WITHIN 0.035 ;
  PROPERTY LEF58_CORNERSPACING "CORNERSPACING CONVEXCORNER EXCEPTEOL 0.08
    WIDTH 0.00 SPACING 0.10
    WIDTH 0.20 SPACING 0.20
    WIDTH 0.50 SPACING 0.30 ;" ;
END Metal7

LAYER Via7
  TYPE CUT ;
  SPACING 0.10 ;
  WIDTH 0.07 ;
  SPACING 0.20 ADJACENTCUTS 3 WITHIN 0.25 ;
END Via7

LAYER Metal8
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.2 0.2 ;
  WIDTH 0.10 ;
  AREA 0.052 ;
  MINWIDTH 0.10 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0.0 0.22 0.47 0.63 1.5
    WIDTH 0	     0.10 0.10 0.10 0.10 0.10
    WIDTH 0.2	     0.10 0.15 0.15 0.15 0.15
    WIDTH 0.4	     0.10 0.15 0.20 0.20 0.20
    WIDTH 1.5	     0.10 0.15 0.20 0.30 0.50 ;
  SPACING 0.12 ENDOFLINE 0.12 WITHIN 0.035 ;
END Metal8

LAYER Via8
  TYPE CUT ;
  SPACING 0.15 ;
  WIDTH 0.10 ;
END Via8

LAYER Metal9
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.2 0.2 ;
  WIDTH 0.10 ;
  AREA 0.052 ;
  MINWIDTH 0.10 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0.0 0.22 0.47 0.63 1.5
    WIDTH 0	     0.10 0.10 0.10 0.10 0.10
    WIDTH 0.2	     0.10 0.15 0.15 0.15 0.15
    WIDTH 0.4	     0.10 0.15 0.20 0.20 0.20
    WIDTH 1.5	     0.10 0.15 0.20 0.30 0.50 ;
  SPACING 0.12 ENDOFLINE 0.12 WITHIN 0.035 ;
END Metal9

LAYER OVERLAP
  TYPE OVERLAP ;
END OVERLAP

VIA VIA12_1C DEFAULT 
    LAYER Metal1 ;
        RECT -0.025000 -0.055000 0.025000 0.055000 ;
    LAYER Via1 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal2 ;
        RECT -0.055000 -0.025000 0.055000 0.025000 ;
END VIA12_1C

VIA VIA12_1C_H DEFAULT 
    LAYER Metal1 ;
        RECT -0.055000 -0.025000 0.055000 0.025000 ;
    LAYER Via1 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal2 ;
        RECT -0.055000 -0.025000 0.055000 0.025000 ;
END VIA12_1C_H

VIA VIA12_1C_V DEFAULT 
    LAYER Metal1 ;
        RECT -0.025000 -0.055000 0.025000 0.055000 ;
    LAYER Via1 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal2 ;
        RECT -0.025000 -0.055000 0.025000 0.055000 ;
END VIA12_1C_V

VIA VIA12_PG
    LAYER Metal1 ;
        RECT -0.350000 -0.050000 0.350000 0.050000 ;
    LAYER Via1 ;
        RECT -0.325000 -0.025000 -0.275000 0.025000 ;
        RECT -0.175000 -0.025000 -0.125000 0.025000 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
        RECT 0.125000 -0.025000 0.175000 0.025000 ;
        RECT 0.275000 -0.025000 0.325000 0.025000 ;
    LAYER Metal2 ;
        RECT -0.350000 -0.050000 0.350000 0.050000 ;
END VIA12_PG

VIA VIA23_1C DEFAULT 
    LAYER Metal2 ;
        RECT -0.055000 -0.025000 0.055000 0.025000 ;
    LAYER Via2 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal3 ;
        RECT -0.025000 -0.055000 0.025000 0.055000 ;
END VIA23_1C

VIA VIA23_1C_H DEFAULT 
    LAYER Metal2 ;
        RECT -0.055000 -0.025000 0.055000 0.025000 ;
    LAYER Via2 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal3 ;
        RECT -0.055000 -0.025000 0.055000 0.025000 ;
END VIA23_1C_H

VIA VIA23_1C_V DEFAULT 
    LAYER Metal2 ;
        RECT -0.025000 -0.055000 0.025000 0.055000 ;
    LAYER Via2 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal3 ;
        RECT -0.025000 -0.055000 0.025000 0.055000 ;
END VIA23_1C_V

VIA VIA23_1ST_E DEFAULT 
    LAYER Metal2 ;
        RECT -0.055000 -0.025000 0.325000 0.025000 ;
    LAYER Via2 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal3 ;
        RECT -0.025000 -0.055000 0.025000 0.055000 ;
END VIA23_1ST_E

VIA VIA23_1ST_W DEFAULT 
    LAYER Metal2 ;
        RECT -0.325000 -0.025000 0.055000 0.025000 ;
    LAYER Via2 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal3 ;
        RECT -0.025000 -0.055000 0.025000 0.055000 ;
END VIA23_1ST_W

VIA VIA23_PG
    LAYER Metal2 ;
        RECT -0.350000 -0.050000 0.350000 0.050000 ;
    LAYER Via2 ;
        RECT -0.325000 -0.025000 -0.275000 0.025000 ;
        RECT -0.175000 -0.025000 -0.125000 0.025000 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
        RECT 0.125000 -0.025000 0.175000 0.025000 ;
        RECT 0.275000 -0.025000 0.325000 0.025000 ;
    LAYER Metal3 ;
        RECT -0.350000 -0.050000 0.350000 0.050000 ;
END VIA23_PG

VIA VIA34_1C DEFAULT 
    LAYER Metal3 ;
        RECT -0.025000 -0.055000 0.025000 0.055000 ;
    LAYER Via3 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal4 ;
        RECT -0.055000 -0.025000 0.055000 0.025000 ;
END VIA34_1C

VIA VIA34_1C_H DEFAULT 
    LAYER Metal3 ;
        RECT -0.055000 -0.025000 0.055000 0.025000 ;
    LAYER Via3 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal4 ;
        RECT -0.055000 -0.025000 0.055000 0.025000 ;
END VIA34_1C_H

VIA VIA34_1C_V DEFAULT 
    LAYER Metal3 ;
        RECT -0.025000 -0.055000 0.025000 0.055000 ;
    LAYER Via3 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal4 ;
        RECT -0.025000 -0.055000 0.025000 0.055000 ;
END VIA34_1C_V

VIA VIA34_1ST_N DEFAULT 
    LAYER Metal3 ;
        RECT -0.025000 -0.055000 0.025000 0.325000 ;
    LAYER Via3 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal4 ;
        RECT -0.055000 -0.025000 0.055000 0.025000 ;
END VIA34_1ST_N

VIA VIA34_1ST_S DEFAULT 
    LAYER Metal3 ;
        RECT -0.025000 -0.325000 0.025000 0.055000 ;
    LAYER Via3 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal4 ;
        RECT -0.055000 -0.025000 0.055000 0.025000 ;
END VIA34_1ST_S

VIA VIA34_PG
    LAYER Metal3 ;
        RECT -0.350000 -0.050000 0.350000 0.050000 ;
    LAYER Via3 ;
        RECT -0.325000 -0.025000 -0.275000 0.025000 ;
        RECT -0.175000 -0.025000 -0.125000 0.025000 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
        RECT 0.125000 -0.025000 0.175000 0.025000 ;
        RECT 0.275000 -0.025000 0.325000 0.025000 ;
    LAYER Metal4 ;
        RECT -0.350000 -0.050000 0.350000 0.050000 ;
END VIA34_PG

VIA VIA45_1C DEFAULT 
    LAYER Metal4 ;
        RECT -0.055000 -0.025000 0.055000 0.025000 ;
    LAYER Via4 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal5 ;
        RECT -0.025000 -0.055000 0.025000 0.055000 ;
END VIA45_1C

VIA VIA45_PG
    LAYER Metal4 ;
        RECT -0.200000 -0.050000 0.200000 0.050000 ;
    LAYER Via4 ;
        RECT -0.175000 -0.025000 -0.125000 0.025000 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
        RECT 0.125000 -0.025000 0.175000 0.025000 ;
    LAYER Metal5 ;
        RECT -0.200000 -0.050000 0.200000 0.050000 ;
END VIA45_PG

VIA VIA5_0_VH DEFAULT 
    LAYER Metal5 ;
        RECT -0.035000 -0.065000 0.035000 0.065000 ;
    LAYER Via5 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal6 ;
        RECT -0.065000 -0.035000 0.065000 0.035000 ;
END VIA5_0_VH

VIA VIA56_PG
    LAYER Metal5 ;
        RECT -0.150000 -0.150000 0.150000 0.150000 ;
    LAYER Via5 ;
        RECT -0.150000 -0.150000 -0.100000 -0.100000 ;
        RECT -0.150000 0.100000 -0.100000 0.150000 ;
        RECT 0.100000 0.100000 0.150000 0.150000 ;
        RECT 0.100000 -0.150000 0.150000 -0.100000 ;
    LAYER Metal6 ;
        RECT -0.150000 -0.150000 0.150000 0.150000 ;
END VIA56_PG

VIA VIA6_0_HV DEFAULT 
    LAYER Metal6 ;
        RECT -0.065000 -0.035000 0.065000 0.035000 ;
    LAYER Via6 ;
        RECT -0.035000 -0.035000 0.035000 0.035000 ;
    LAYER Metal7 ;
        RECT -0.035000 -0.065000 0.035000 0.065000 ;
END VIA6_0_HV

VIA VIA67_PG
    LAYER Metal6 ;
        RECT -0.170000 -0.170000 0.170000 0.170000 ;
    LAYER Via6 ;
        RECT -0.170000 -0.170000 -0.100000 -0.100000 ;
        RECT -0.170000 0.100000 -0.100000 0.170000 ;
        RECT 0.100000 0.100000 0.170000 0.170000 ;
        RECT 0.100000 -0.170000 0.170000 -0.100000 ;
    LAYER Metal7 ;
        RECT -0.170000 -0.170000 0.170000 0.170000 ;
END VIA67_PG

VIA VIA7_0_VH DEFAULT 
    LAYER Metal7 ;
        RECT -0.050000 -0.260000 0.050000 0.260000 ;
    LAYER Via7 ;
        RECT -0.050000 -0.050000 0.050000 0.050000 ;
    LAYER Metal8 ;
        RECT -0.260000 -0.050000 0.260000 0.050000 ;
END VIA7_0_VH

VIA VIA78_PG
    LAYER Metal7 ;
        RECT -0.170000 -0.170000 0.170000 0.170000 ;
    LAYER Via7 ;
        RECT -0.170000 -0.170000 -0.100000 -0.100000 ;
        RECT -0.170000 0.100000 -0.100000 0.170000 ;
        RECT 0.100000 0.100000 0.170000 0.170000 ;
        RECT 0.100000 -0.170000 0.170000 -0.100000 ;
    LAYER Metal8 ;
        RECT -0.170000 -0.170000 0.170000 0.170000 ;
END VIA78_PG

VIA VIA8_0_HV DEFAULT 
    LAYER Metal8 ;
        RECT -0.260000 -0.050000 0.260000 0.050000 ;
    LAYER Via8 ;
        RECT -0.050000 -0.050000 0.050000 0.050000 ;
    LAYER Metal9 ;
        RECT -0.050000 -0.260000 0.050000 0.260000 ;
END VIA8_0_HV

SITE CoreSite
  CLASS CORE ;
  SIZE 0.1 BY 1.2 ;
END CoreSite


MACRO XOR2X1
    CLASS CORE ;
    FOREIGN XOR2X1 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.400000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.440000 0.557000 0.542000 0.638000 ;
        RECT 0.162000 0.433000 0.232000 0.496000 ;
        RECT 0.440000 0.439000 0.501000 0.638000 ;
        RECT 0.162000 0.388000 0.223000 0.496000 ;
        RECT 0.407000 0.439000 0.501000 0.496000 ;
        RECT 0.162000 0.442000 0.501000 0.496000 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.289000 0.570000 0.350000 0.761000 ;
        RECT 0.289000 0.570000 0.379000 0.625000 ;
        RECT 0.232000 0.706000 0.350000 0.761000 ;
        END
    END B
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 1.400000 1.280000 ;
        RECT 1.114000 1.078000 1.204000 1.280000 ;
        RECT 0.215000 1.078000 0.305000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 1.400000 0.080000 ;
        RECT 1.114000 -0.080000 1.204000 0.122000 ;
        RECT 0.235000 -0.080000 0.325000 0.122000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.262000 0.707000 1.352000 0.788000 ;
        RECT 1.262000 0.279000 1.352000 0.360000 ;
        RECT 1.282000 0.573000 1.352000 0.788000 ;
        RECT 1.291000 0.279000 1.352000 0.788000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.040000 0.810000 0.138000 0.901000 ;
        RECT 0.973000 0.858000 1.063000 0.974000 ;
        RECT 0.927000 0.702000 1.035000 0.789000 ;
        RECT 1.126000 0.426000 1.229000 0.507000 ;
        RECT 0.477000 0.745000 0.664000 0.826000 ;
        RECT 1.126000 0.194000 1.187000 0.507000 ;
        RECT 0.974000 0.304000 1.035000 0.789000 ;
        RECT 0.736000 0.194000 0.797000 0.802000 ;
        RECT 0.603000 0.311000 0.664000 0.913000 ;
        RECT 0.386000 0.150000 0.447000 0.246000 ;
        RECT 0.366000 0.902000 0.427000 1.029000 ;
        RECT 0.077000 0.810000 0.138000 0.957000 ;
        RECT 0.077000 0.192000 0.138000 0.313000 ;
        RECT 0.040000 0.258000 0.101000 0.901000 ;
        RECT 0.736000 0.194000 1.187000 0.249000 ;
        RECT 0.603000 0.858000 1.063000 0.913000 ;
        RECT 0.386000 0.150000 0.675000 0.205000 ;
        RECT 0.366000 0.974000 0.875000 1.029000 ;
        RECT 0.077000 0.902000 0.427000 0.957000 ;
        RECT 0.040000 0.258000 0.138000 0.313000 ;
        RECT 0.912000 0.304000 1.035000 0.358000 ;
        RECT 0.477000 0.311000 0.664000 0.365000 ;
        RECT 0.077000 0.192000 0.447000 0.246000 ;
        RECT 0.077000 0.192000 0.101000 0.957000 ;
    END
END XOR2X1

MACRO SEDFFHQX2
    CLASS CORE ;
    FOREIGN SEDFFHQX2 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 5.900000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER Metal1 ;
        RECT 2.448000 0.421000 2.628000 0.512000 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.078000 0.433000 1.179000 0.564000 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.772000 0.549000 1.872000 0.693000 ;
        RECT 1.702000 0.555000 1.872000 0.610000 ;
        END
    END E
    PIN Q
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 5.763000 0.652000 5.862000 0.767000 ;
        RECT 5.758000 0.652000 5.863000 0.733000 ;
        RECT 5.758000 0.346000 5.863000 0.427000 ;
        RECT 5.803000 0.346000 5.863000 0.733000 ;
        RECT 5.803000 0.346000 5.862000 0.767000 ;
        END
    END Q
    PIN SE
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.170000 0.490000 0.291000 0.633000 ;
        END
    END SE
    PIN SI
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.371000 0.167000 0.511000 0.262000 ;
        END
    END SI
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 5.900000 1.280000 ;
        RECT 5.579000 1.078000 5.669000 1.280000 ;
        RECT 5.186000 1.078000 5.276000 1.280000 ;
        RECT 1.727000 1.078000 1.817000 1.280000 ;
        RECT 1.021000 1.078000 1.111000 1.280000 ;
        RECT 3.149000 1.078000 3.238000 1.280000 ;
        RECT 0.221000 1.078000 0.310000 1.280000 ;
        RECT 2.624000 0.902000 2.684000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 5.900000 0.080000 ;
        RECT 5.579000 -0.080000 5.669000 0.122000 ;
        RECT 3.340000 -0.080000 3.430000 0.287000 ;
        RECT 1.731000 -0.080000 1.821000 0.122000 ;
        RECT 5.205000 -0.080000 5.294000 0.122000 ;
        RECT 4.311000 -0.080000 4.400000 0.395000 ;
        RECT 3.932000 -0.080000 4.021000 0.342000 ;
        RECT 2.641000 -0.080000 2.730000 0.122000 ;
        RECT 1.024000 -0.080000 1.113000 0.122000 ;
        RECT 0.205000 -0.080000 0.294000 0.122000 ;
        END
    END VSS
    OBS
        LAYER Metal1 ;
        RECT 5.404000 0.748000 5.494000 0.940000 ;
        RECT 1.956000 0.542000 2.068000 0.631000 ;
        RECT 1.520000 0.526000 1.612000 0.613000 ;
        RECT 0.785000 0.469000 0.885000 0.554000 ;
        RECT 5.652000 0.500000 5.741000 0.581000 ;
        RECT 5.404000 0.292000 5.494000 0.373000 ;
        RECT 5.278000 0.543000 5.368000 0.624000 ;
        RECT 4.121000 0.276000 4.211000 0.357000 ;
        RECT 2.983000 0.255000 3.072000 0.336000 ;
        RECT 2.436000 0.231000 2.525000 0.312000 ;
        RECT 1.942000 0.668000 2.031000 0.749000 ;
        RECT 1.566000 0.668000 1.655000 0.749000 ;
        RECT 1.361000 0.287000 1.450000 0.368000 ;
        RECT 1.171000 0.657000 1.261000 0.738000 ;
        RECT 1.171000 0.287000 1.261000 0.368000 ;
        RECT 0.626000 0.343000 0.715000 0.424000 ;
        RECT 0.594000 0.820000 0.684000 0.901000 ;
        RECT 0.455000 0.969000 0.544000 1.050000 ;
        RECT 0.415000 0.343000 0.505000 0.424000 ;
        RECT 0.394000 0.746000 0.484000 0.827000 ;
        RECT 0.047000 0.343000 0.137000 0.424000 ;
        RECT 5.278000 0.543000 5.353000 0.627000 ;
        RECT 4.852000 0.814000 4.927000 0.927000 ;
        RECT 1.956000 0.542000 2.031000 0.749000 ;
        RECT 0.455000 0.935000 0.530000 1.050000 ;
        RECT 2.063000 0.833000 2.190000 0.902000 ;
        RECT 5.432000 0.526000 5.494000 0.940000 ;
        RECT 5.116000 0.683000 5.177000 0.910000 ;
        RECT 5.053000 0.855000 5.114000 1.050000 ;
        RECT 5.031000 0.174000 5.092000 0.268000 ;
        RECT 4.973000 0.573000 5.034000 0.773000 ;
        RECT 4.881000 0.718000 4.942000 0.895000 ;
        RECT 4.840000 0.330000 4.901000 0.649000 ;
        RECT 4.609000 0.261000 4.670000 0.792000 ;
        RECT 4.488000 0.735000 4.549000 0.927000 ;
        RECT 4.472000 0.150000 4.533000 0.242000 ;
        RECT 4.338000 0.594000 4.399000 0.940000 ;
        RECT 3.544000 0.231000 3.605000 0.831000 ;
        RECT 3.030000 0.268000 3.091000 0.650000 ;
        RECT 2.266000 0.306000 2.327000 0.915000 ;
        RECT 2.077000 0.306000 2.138000 0.445000 ;
        RECT 1.956000 0.150000 2.017000 0.749000 ;
        RECT 1.911000 0.954000 1.972000 1.037000 ;
        RECT 1.551000 0.302000 1.612000 0.736000 ;
        RECT 1.551000 0.161000 1.612000 0.246000 ;
        RECT 1.375000 0.287000 1.436000 0.899000 ;
        RECT 0.828000 0.163000 0.889000 0.257000 ;
        RECT 0.824000 0.318000 0.885000 0.733000 ;
        RECT 0.623000 0.820000 0.684000 1.008000 ;
        RECT 0.415000 0.343000 0.476000 0.827000 ;
        RECT 0.076000 0.746000 0.137000 0.989000 ;
        RECT 0.047000 0.343000 0.108000 0.827000 ;
        RECT 5.432000 0.292000 5.492000 0.940000 ;
        RECT 5.105000 0.213000 5.165000 0.627000 ;
        RECT 4.834000 0.150000 4.894000 0.229000 ;
        RECT 4.136000 0.276000 4.196000 0.805000 ;
        RECT 4.010000 0.508000 4.070000 0.831000 ;
        RECT 3.681000 0.289000 3.741000 0.720000 ;
        RECT 3.422000 0.843000 3.482000 0.940000 ;
        RECT 3.418000 0.357000 3.478000 0.462000 ;
        RECT 3.300000 0.954000 3.360000 1.050000 ;
        RECT 2.987000 0.595000 3.047000 0.783000 ;
        RECT 2.866000 0.665000 2.926000 0.898000 ;
        RECT 2.745000 0.776000 2.805000 1.008000 ;
        RECT 2.698000 0.257000 2.758000 0.720000 ;
        RECT 2.130000 0.390000 2.190000 0.902000 ;
        RECT 1.830000 0.375000 1.890000 0.482000 ;
        RECT 1.240000 0.300000 1.300000 0.725000 ;
        RECT 0.947000 0.202000 1.007000 0.899000 ;
        RECT 0.626000 0.343000 0.686000 0.501000 ;
        RECT 0.609000 0.446000 0.669000 0.901000 ;
        RECT 5.432000 0.526000 5.741000 0.581000 ;
        RECT 5.053000 0.855000 5.494000 0.910000 ;
        RECT 5.031000 0.213000 5.165000 0.268000 ;
        RECT 4.881000 0.718000 5.034000 0.773000 ;
        RECT 4.840000 0.330000 5.038000 0.385000 ;
        RECT 4.834000 0.174000 5.092000 0.229000 ;
        RECT 4.730000 0.594000 4.901000 0.649000 ;
        RECT 4.609000 0.737000 4.752000 0.792000 ;
        RECT 4.472000 0.150000 4.894000 0.205000 ;
        RECT 4.338000 0.594000 4.545000 0.649000 ;
        RECT 4.136000 0.470000 4.670000 0.525000 ;
        RECT 3.681000 0.665000 3.832000 0.720000 ;
        RECT 3.681000 0.289000 3.832000 0.344000 ;
        RECT 3.544000 0.776000 4.070000 0.831000 ;
        RECT 3.300000 0.995000 5.114000 1.050000 ;
        RECT 3.030000 0.357000 3.478000 0.412000 ;
        RECT 2.866000 0.843000 3.482000 0.898000 ;
        RECT 2.698000 0.394000 2.964000 0.449000 ;
        RECT 2.436000 0.257000 2.758000 0.312000 ;
        RECT 2.410000 0.665000 2.926000 0.720000 ;
        RECT 2.266000 0.776000 2.805000 0.831000 ;
        RECT 1.956000 0.150000 2.052000 0.205000 ;
        RECT 1.911000 0.982000 2.440000 1.037000 ;
        RECT 1.551000 0.427000 1.890000 0.482000 ;
        RECT 1.551000 0.302000 1.647000 0.357000 ;
        RECT 1.375000 0.833000 2.190000 0.888000 ;
        RECT 0.828000 0.202000 1.007000 0.257000 ;
        RECT 0.797000 0.844000 1.436000 0.899000 ;
        RECT 0.797000 0.163000 0.889000 0.218000 ;
        RECT 4.973000 0.573000 5.353000 0.627000 ;
        RECT 4.609000 0.261000 4.737000 0.315000 ;
        RECT 4.488000 0.873000 4.927000 0.927000 ;
        RECT 3.422000 0.886000 4.399000 0.940000 ;
        RECT 3.233000 0.554000 3.605000 0.608000 ;
        RECT 2.745000 0.954000 3.360000 1.008000 ;
        RECT 1.551000 0.192000 2.017000 0.246000 ;
        RECT 1.298000 0.161000 1.612000 0.215000 ;
        RECT 0.623000 0.954000 1.972000 1.008000 ;
        RECT 0.076000 0.935000 0.530000 0.989000 ;
        RECT 4.881000 0.718000 4.927000 0.927000 ;
        RECT 1.566000 0.302000 1.612000 0.749000 ;
        RECT 0.623000 0.446000 0.669000 1.008000 ;
        RECT 0.626000 0.343000 0.669000 1.008000 ;
        RECT 3.030000 0.255000 3.072000 0.650000 ;
        RECT 0.076000 0.343000 0.108000 0.989000 ;
        RECT 1.240000 0.287000 1.261000 0.738000 ;
        RECT 3.030000 0.255000 3.047000 0.783000 ;
        RECT 2.130000 0.306000 2.138000 0.902000 ;
    END
END SEDFFHQX2

MACRO SEDFFHQX1
    CLASS CORE ;
    FOREIGN SEDFFHQX1 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 5.400000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER Metal1 ;
        RECT 2.457000 0.421000 2.638000 0.512000 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.082000 0.433000 1.184000 0.564000 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.779000 0.549000 1.879000 0.693000 ;
        RECT 1.709000 0.555000 1.879000 0.610000 ;
        END
    END E
    PIN Q
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 5.251000 0.690000 5.343000 0.771000 ;
        RECT 5.227000 0.324000 5.343000 0.405000 ;
        RECT 5.283000 0.324000 5.343000 0.771000 ;
        END
    END Q
    PIN SE
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.170000 0.490000 0.292000 0.633000 ;
        END
    END SE
    PIN SI
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.372000 0.167000 0.513000 0.262000 ;
        END
    END SI
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 5.400000 1.280000 ;
        RECT 5.081000 1.078000 5.194000 1.280000 ;
        RECT 4.716000 1.078000 4.806000 1.280000 ;
        RECT 1.734000 1.078000 1.824000 1.280000 ;
        RECT 1.025000 1.078000 1.115000 1.280000 ;
        RECT 3.161000 1.078000 3.250000 1.280000 ;
        RECT 0.222000 1.078000 0.311000 1.280000 ;
        RECT 2.634000 0.902000 2.695000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 5.400000 0.080000 ;
        RECT 5.079000 -0.080000 5.169000 0.122000 ;
        RECT 4.727000 -0.080000 4.817000 0.122000 ;
        RECT 3.947000 -0.080000 4.037000 0.370000 ;
        RECT 3.332000 -0.080000 3.422000 0.287000 ;
        RECT 2.651000 -0.080000 2.741000 0.122000 ;
        RECT 1.738000 -0.080000 1.828000 0.122000 ;
        RECT 1.028000 -0.080000 1.118000 0.122000 ;
        RECT 0.206000 -0.080000 0.296000 0.122000 ;
        END
    END VSS
    OBS
        LAYER Metal1 ;
        RECT 4.918000 0.742000 5.008000 0.935000 ;
        RECT 1.964000 0.542000 2.076000 0.631000 ;
        RECT 1.526000 0.526000 1.618000 0.613000 ;
        RECT 0.788000 0.469000 0.888000 0.554000 ;
        RECT 5.124000 0.500000 5.214000 0.581000 ;
        RECT 4.895000 0.307000 4.984000 0.388000 ;
        RECT 4.757000 0.524000 4.847000 0.605000 ;
        RECT 4.632000 0.683000 4.722000 0.764000 ;
        RECT 2.445000 0.231000 2.535000 0.312000 ;
        RECT 0.417000 0.343000 0.507000 0.424000 ;
        RECT 0.396000 0.746000 0.486000 0.827000 ;
        RECT 0.048000 0.746000 0.137000 0.827000 ;
        RECT 0.048000 0.343000 0.137000 0.424000 ;
        RECT 4.603000 0.480000 4.679000 0.579000 ;
        RECT 4.924000 0.513000 4.994000 0.935000 ;
        RECT 2.071000 0.833000 2.199000 0.902000 ;
        RECT 4.646000 0.683000 4.707000 0.910000 ;
        RECT 4.603000 0.151000 4.664000 0.579000 ;
        RECT 4.394000 0.855000 4.455000 1.050000 ;
        RECT 4.394000 0.717000 4.455000 0.800000 ;
        RECT 4.278000 0.332000 4.339000 0.669000 ;
        RECT 4.273000 0.614000 4.334000 0.940000 ;
        RECT 4.025000 0.508000 4.086000 0.831000 ;
        RECT 3.699000 0.150000 3.760000 0.720000 ;
        RECT 3.435000 0.843000 3.496000 0.940000 ;
        RECT 3.431000 0.357000 3.492000 0.462000 ;
        RECT 3.312000 0.954000 3.373000 1.050000 ;
        RECT 2.998000 0.595000 3.059000 0.783000 ;
        RECT 2.877000 0.665000 2.938000 0.898000 ;
        RECT 2.755000 0.776000 2.816000 1.008000 ;
        RECT 2.275000 0.306000 2.336000 0.915000 ;
        RECT 2.138000 0.390000 2.199000 0.902000 ;
        RECT 2.085000 0.306000 2.146000 0.445000 ;
        RECT 1.837000 0.375000 1.898000 0.482000 ;
        RECT 1.557000 0.302000 1.618000 0.736000 ;
        RECT 1.557000 0.161000 1.618000 0.246000 ;
        RECT 1.380000 0.287000 1.441000 0.888000 ;
        RECT 0.950000 0.202000 1.011000 0.888000 ;
        RECT 0.831000 0.163000 0.892000 0.257000 ;
        RECT 0.827000 0.318000 0.888000 0.733000 ;
        RECT 0.611000 0.446000 0.672000 1.008000 ;
        RECT 0.471000 0.935000 0.532000 1.050000 ;
        RECT 0.417000 0.343000 0.478000 0.827000 ;
        RECT 4.924000 0.307000 4.984000 0.935000 ;
        RECT 4.482000 0.298000 4.542000 0.387000 ;
        RECT 4.404000 0.480000 4.464000 0.771000 ;
        RECT 4.342000 0.151000 4.402000 0.268000 ;
        RECT 4.152000 0.271000 4.212000 0.780000 ;
        RECT 3.558000 0.233000 3.618000 0.831000 ;
        RECT 3.042000 0.244000 3.102000 0.650000 ;
        RECT 2.699000 0.257000 2.759000 0.720000 ;
        RECT 1.964000 0.150000 2.024000 0.749000 ;
        RECT 1.919000 0.954000 1.979000 1.037000 ;
        RECT 1.246000 0.300000 1.306000 0.725000 ;
        RECT 0.643000 0.343000 0.703000 0.501000 ;
        RECT 0.077000 0.746000 0.137000 0.989000 ;
        RECT 0.048000 0.343000 0.108000 0.827000 ;
        RECT 4.278000 0.332000 4.334000 0.940000 ;
        RECT 4.994000 0.513000 5.214000 0.568000 ;
        RECT 4.924000 0.513000 5.008000 0.568000 ;
        RECT 4.603000 0.524000 4.847000 0.579000 ;
        RECT 4.404000 0.480000 4.679000 0.535000 ;
        RECT 4.394000 0.855000 5.008000 0.910000 ;
        RECT 4.342000 0.151000 4.664000 0.206000 ;
        RECT 4.278000 0.332000 4.542000 0.387000 ;
        RECT 4.273000 0.614000 4.339000 0.669000 ;
        RECT 3.699000 0.665000 3.847000 0.720000 ;
        RECT 3.558000 0.776000 4.086000 0.831000 ;
        RECT 3.312000 0.995000 4.455000 1.050000 ;
        RECT 3.245000 0.357000 3.492000 0.412000 ;
        RECT 3.102000 0.357000 3.431000 0.412000 ;
        RECT 3.042000 0.357000 3.373000 0.412000 ;
        RECT 2.998000 0.595000 3.102000 0.650000 ;
        RECT 2.973000 0.244000 3.102000 0.299000 ;
        RECT 2.877000 0.843000 3.496000 0.898000 ;
        RECT 2.699000 0.394000 2.965000 0.449000 ;
        RECT 2.445000 0.257000 2.759000 0.312000 ;
        RECT 2.419000 0.776000 2.816000 0.831000 ;
        RECT 2.419000 0.665000 2.938000 0.720000 ;
        RECT 2.336000 0.776000 2.755000 0.831000 ;
        RECT 2.275000 0.776000 2.699000 0.831000 ;
        RECT 2.085000 0.390000 2.199000 0.445000 ;
        RECT 1.964000 0.150000 2.060000 0.205000 ;
        RECT 1.919000 0.982000 2.449000 1.037000 ;
        RECT 1.557000 0.681000 1.661000 0.736000 ;
        RECT 1.557000 0.427000 1.898000 0.482000 ;
        RECT 1.557000 0.302000 1.654000 0.357000 ;
        RECT 1.176000 0.670000 1.306000 0.725000 ;
        RECT 1.176000 0.300000 1.306000 0.355000 ;
        RECT 0.831000 0.202000 1.011000 0.257000 ;
        RECT 0.800000 0.833000 2.199000 0.888000 ;
        RECT 0.800000 0.163000 0.892000 0.218000 ;
        RECT 0.611000 0.446000 0.703000 0.501000 ;
        RECT 4.394000 0.717000 4.464000 0.771000 ;
        RECT 3.699000 0.317000 3.826000 0.371000 ;
        RECT 3.435000 0.886000 4.334000 0.940000 ;
        RECT 3.245000 0.554000 3.618000 0.608000 ;
        RECT 2.755000 0.954000 3.373000 1.008000 ;
        RECT 1.557000 0.192000 2.024000 0.246000 ;
        RECT 1.302000 0.161000 1.618000 0.215000 ;
        RECT 0.611000 0.954000 1.979000 1.008000 ;
        RECT 0.077000 0.935000 0.532000 0.989000 ;
        RECT 4.404000 0.480000 4.455000 0.800000 ;
        RECT 0.077000 0.343000 0.108000 0.989000 ;
        RECT 0.643000 0.343000 0.672000 1.008000 ;
        RECT 3.042000 0.244000 3.059000 0.783000 ;
        RECT 2.138000 0.306000 2.146000 0.902000 ;
    END
END SEDFFHQX1

MACRO SDFFHQX4
    CLASS CORE ;
    FOREIGN SDFFHQX4 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 4.500000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER Metal1 ;
        RECT 0.152000 0.524000 0.290000 0.627000 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.067000 0.356000 1.156000 0.437000 ;
        RECT 1.088000 0.356000 1.156000 0.439000 ;
        RECT 1.088000 0.356000 1.150000 0.627000 ;
        RECT 1.088000 0.573000 1.155000 0.627000 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 4.191000 0.433000 4.290000 0.767000 ;
        RECT 4.193000 0.325000 4.282000 0.767000 ;
        RECT 4.130000 0.671000 4.290000 0.752000 ;
        END
    END Q
    PIN SE
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.926000 0.593000 1.015000 0.674000 ;
        RECT 0.527000 0.567000 0.690000 0.633000 ;
        RECT 0.629000 0.567000 0.690000 0.656000 ;
        RECT 0.629000 0.601000 1.015000 0.656000 ;
        END
    END SE
    PIN SI
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.750000 0.433000 0.871000 0.533000 ;
        RECT 0.750000 0.433000 0.839000 0.546000 ;
        RECT 0.729000 0.433000 0.871000 0.500000 ;
        END
    END SI
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 3.060000 1.078000 3.687000 1.280000 ;
        RECT 0.000000 1.120000 4.500000 1.280000 ;
        RECT 4.299000 0.989000 4.389000 1.280000 ;
        RECT 3.951000 1.078000 4.040000 1.280000 ;
        RECT 2.284000 1.078000 2.373000 1.280000 ;
        RECT 1.390000 1.078000 1.479000 1.280000 ;
        RECT 0.248000 1.078000 0.337000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 4.500000 0.080000 ;
        RECT 4.025000 -0.080000 4.115000 0.212000 ;
        RECT 4.361000 -0.080000 4.450000 0.215000 ;
        RECT 3.632000 -0.080000 3.721000 0.122000 ;
        RECT 1.678000 -0.080000 1.767000 0.287000 ;
        RECT 0.755000 -0.080000 0.844000 0.122000 ;
        RECT 0.249000 -0.080000 0.338000 0.410000 ;
        RECT 2.361000 -0.080000 2.422000 0.311000 ;
        RECT 3.185000 -0.080000 3.245000 0.287000 ;
        RECT 0.249000 0.359000 0.346000 0.410000 ;
        END
    END VSS
    OBS
        LAYER Metal1 ;
        RECT 0.399000 0.154000 0.490000 0.246000 ;
        RECT 0.490000 0.318000 0.580000 0.425000 ;
        RECT 3.380000 0.150000 3.469000 0.412000 ;
        RECT 2.596000 0.605000 2.685000 0.787000 ;
        RECT 0.047000 0.739000 0.136000 0.932000 ;
        RECT 0.406000 0.692000 0.509000 0.779000 ;
        RECT 1.112000 0.160000 1.201000 0.246000 ;
        RECT 3.842000 0.264000 3.931000 0.345000 ;
        RECT 3.842000 0.264000 3.923000 0.571000 ;
        RECT 3.799000 0.826000 3.923000 0.907000 ;
        RECT 3.699000 0.490000 3.923000 0.571000 ;
        RECT 3.576000 0.650000 3.802000 0.731000 ;
        RECT 3.265000 0.577000 3.354000 0.658000 ;
        RECT 2.913000 0.348000 3.003000 0.429000 ;
        RECT 2.911000 0.596000 3.000000 0.677000 ;
        RECT 2.725000 0.223000 2.814000 0.304000 ;
        RECT 2.672000 0.954000 2.761000 1.035000 ;
        RECT 2.536000 0.245000 2.628000 0.326000 ;
        RECT 2.483000 0.843000 2.573000 0.924000 ;
        RECT 2.420000 0.490000 2.510000 0.571000 ;
        RECT 2.221000 0.504000 2.310000 0.585000 ;
        RECT 2.137000 0.789000 2.226000 0.870000 ;
        RECT 2.010000 0.454000 2.161000 0.535000 ;
        RECT 1.952000 0.790000 2.042000 0.871000 ;
        RECT 1.867000 0.273000 1.956000 0.354000 ;
        RECT 1.740000 0.450000 1.829000 0.531000 ;
        RECT 1.689000 0.612000 1.950000 0.693000 ;
        RECT 1.545000 0.938000 1.634000 1.019000 ;
        RECT 1.248000 0.331000 1.337000 0.412000 ;
        RECT 1.193000 0.776000 1.282000 0.857000 ;
        RECT 0.606000 0.724000 0.695000 0.805000 ;
        RECT 0.068000 0.344000 0.157000 0.425000 ;
        RECT 0.047000 0.688000 0.122000 0.932000 ;
        RECT 1.889000 0.790000 2.042000 0.858000 ;
        RECT 3.414000 0.467000 3.475000 0.768000 ;
        RECT 3.064000 0.223000 3.125000 0.412000 ;
        RECT 3.060000 0.604000 3.121000 0.787000 ;
        RECT 2.942000 0.348000 3.003000 0.521000 ;
        RECT 2.567000 0.245000 2.628000 0.429000 ;
        RECT 2.420000 0.381000 2.481000 0.571000 ;
        RECT 2.137000 0.679000 2.198000 0.870000 ;
        RECT 2.120000 0.269000 2.181000 0.402000 ;
        RECT 1.889000 0.273000 1.950000 0.858000 ;
        RECT 1.463000 0.163000 1.524000 0.855000 ;
        RECT 1.084000 0.939000 1.145000 1.050000 ;
        RECT 0.490000 0.318000 0.551000 0.512000 ;
        RECT 0.422000 0.877000 0.483000 1.050000 ;
        RECT 0.406000 0.457000 0.467000 0.779000 ;
        RECT 0.031000 0.369000 0.092000 0.743000 ;
        RECT 3.863000 0.264000 3.923000 0.907000 ;
        RECT 3.576000 0.357000 3.636000 0.886000 ;
        RECT 3.303000 0.831000 3.363000 1.008000 ;
        RECT 3.181000 0.713000 3.241000 0.898000 ;
        RECT 2.747000 0.490000 2.807000 0.652000 ;
        RECT 2.287000 0.530000 2.347000 0.993000 ;
        RECT 2.241000 0.158000 2.301000 0.436000 ;
        RECT 2.101000 0.348000 2.161000 0.733000 ;
        RECT 1.896000 0.158000 1.956000 0.354000 ;
        RECT 1.343000 0.357000 1.403000 0.994000 ;
        RECT 0.952000 0.802000 1.012000 0.936000 ;
        RECT 0.031000 0.369000 0.157000 0.425000 ;
        RECT 3.303000 0.831000 3.636000 0.886000 ;
        RECT 3.181000 0.713000 3.475000 0.768000 ;
        RECT 3.064000 0.357000 3.636000 0.412000 ;
        RECT 2.567000 0.374000 3.003000 0.429000 ;
        RECT 2.483000 0.843000 3.241000 0.898000 ;
        RECT 2.483000 0.490000 2.807000 0.545000 ;
        RECT 2.420000 0.490000 2.725000 0.545000 ;
        RECT 2.287000 0.732000 3.121000 0.787000 ;
        RECT 2.241000 0.381000 2.481000 0.436000 ;
        RECT 2.221000 0.530000 2.347000 0.585000 ;
        RECT 1.896000 0.158000 2.301000 0.213000 ;
        RECT 1.545000 0.938000 2.347000 0.993000 ;
        RECT 1.545000 0.450000 1.829000 0.505000 ;
        RECT 1.524000 0.450000 1.740000 0.505000 ;
        RECT 1.463000 0.450000 1.689000 0.505000 ;
        RECT 1.322000 0.163000 1.524000 0.218000 ;
        RECT 1.248000 0.357000 1.403000 0.412000 ;
        RECT 1.084000 0.939000 1.634000 0.994000 ;
        RECT 0.952000 0.802000 1.282000 0.857000 ;
        RECT 0.543000 0.881000 1.012000 0.936000 ;
        RECT 0.490000 0.318000 0.952000 0.373000 ;
        RECT 0.422000 0.995000 1.145000 1.050000 ;
        RECT 0.406000 0.724000 0.695000 0.779000 ;
        RECT 0.406000 0.457000 0.551000 0.512000 ;
        RECT 0.047000 0.877000 0.483000 0.932000 ;
        RECT 0.031000 0.688000 0.122000 0.743000 ;
        RECT 3.060000 0.604000 3.354000 0.658000 ;
        RECT 2.942000 0.467000 3.475000 0.521000 ;
        RECT 2.747000 0.598000 3.000000 0.652000 ;
        RECT 2.725000 0.223000 3.125000 0.277000 ;
        RECT 2.672000 0.954000 3.363000 1.008000 ;
        RECT 2.101000 0.679000 2.198000 0.733000 ;
        RECT 2.101000 0.348000 2.181000 0.402000 ;
        RECT 1.896000 0.158000 1.950000 0.858000 ;
        RECT 1.084000 0.939000 2.347000 0.993000 ;
        RECT 0.399000 0.192000 1.201000 0.246000 ;
        RECT 2.137000 0.269000 2.161000 0.870000 ;
        RECT 0.068000 0.344000 0.092000 0.932000 ;
        RECT 2.287000 0.504000 2.310000 0.993000 ;
        RECT 0.047000 0.369000 0.068000 0.932000 ;
        RECT 2.120000 0.269000 2.137000 0.733000 ;
    END
END SDFFHQX4

MACRO SDFFHQX2
    CLASS CORE ;
    FOREIGN SDFFHQX2 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 4.200000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER Metal1 ;
        RECT 0.212000 0.512000 0.327000 0.633000 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.051000 0.335000 1.184000 0.494000 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 3.855000 0.167000 3.945000 0.248000 ;
        RECT 3.695000 0.700000 3.813000 0.767000 ;
        RECT 3.695000 0.193000 3.756000 0.767000 ;
        RECT 3.695000 0.193000 3.945000 0.248000 ;
        END
    END Q
    PIN SE
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.998000 0.648000 1.088000 0.729000 ;
        RECT 0.562000 0.567000 0.663000 0.635000 ;
        RECT 0.544000 0.568000 0.663000 0.635000 ;
        RECT 0.998000 0.574000 1.059000 0.729000 ;
        RECT 0.544000 0.574000 1.059000 0.629000 ;
        END
    END SE
    PIN SI
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.655000 0.412000 0.790000 0.500000 ;
        RECT 0.655000 0.433000 0.838000 0.500000 ;
        END
    END SI
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 2.983000 1.078000 3.447000 1.280000 ;
        RECT 0.000000 1.120000 4.200000 1.280000 ;
        RECT 3.882000 1.078000 3.972000 1.280000 ;
        RECT 2.182000 1.078000 2.272000 1.280000 ;
        RECT 0.997000 1.065000 1.087000 1.280000 ;
        RECT 0.313000 1.078000 0.403000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 4.200000 0.080000 ;
        RECT 0.742000 -0.080000 0.833000 0.122000 ;
        RECT 4.057000 -0.080000 4.147000 0.211000 ;
        RECT 3.643000 -0.080000 3.733000 0.122000 ;
        RECT 2.286000 -0.080000 2.376000 0.308000 ;
        RECT 1.676000 -0.080000 1.766000 0.287000 ;
        RECT 0.231000 -0.080000 0.321000 0.409000 ;
        RECT 3.138000 -0.080000 3.199000 0.241000 ;
        RECT 0.231000 0.358000 0.329000 0.409000 ;
        END
    END VSS
    OBS
        LAYER Metal1 ;
        RECT 0.103000 0.719000 0.209000 0.913000 ;
        RECT 3.679000 0.931000 3.770000 1.040000 ;
        RECT 3.336000 0.277000 3.426000 0.412000 ;
        RECT 2.591000 0.576000 2.681000 0.752000 ;
        RECT 1.588000 0.926000 1.677000 1.019000 ;
        RECT 2.039000 0.150000 2.125000 0.344000 ;
        RECT 1.588000 0.933000 1.678000 1.019000 ;
        RECT 3.855000 0.348000 3.945000 0.429000 ;
        RECT 3.367000 0.917000 3.458000 0.998000 ;
        RECT 3.116000 0.800000 3.206000 0.881000 ;
        RECT 2.781000 0.807000 2.872000 0.888000 ;
        RECT 2.591000 0.917000 2.681000 0.998000 ;
        RECT 2.487000 0.262000 2.577000 0.343000 ;
        RECT 2.039000 0.263000 2.164000 0.344000 ;
        RECT 1.661000 0.514000 1.963000 0.595000 ;
        RECT 1.315000 0.193000 1.405000 0.274000 ;
        RECT 1.266000 0.769000 1.356000 0.850000 ;
        RECT 1.254000 0.329000 1.344000 0.410000 ;
        RECT 1.103000 0.179000 1.193000 0.260000 ;
        RECT 0.602000 0.724000 0.692000 0.805000 ;
        RECT 0.472000 0.343000 0.562000 0.424000 ;
        RECT 0.048000 0.319000 0.151000 0.400000 ;
        RECT 0.419000 0.700000 0.552000 0.779000 ;
        RECT 0.487000 0.302000 0.562000 0.424000 ;
        RECT 0.851000 0.302000 0.941000 0.373000 ;
        RECT 0.090000 0.719000 0.209000 0.788000 ;
        RECT 1.417000 0.926000 1.677000 0.988000 ;
        RECT 3.997000 0.374000 4.058000 0.986000 ;
        RECT 3.874000 0.544000 3.935000 0.876000 ;
        RECT 3.573000 0.357000 3.634000 0.876000 ;
        RECT 3.451000 0.467000 3.512000 0.745000 ;
        RECT 3.116000 0.800000 3.177000 0.998000 ;
        RECT 3.005000 0.152000 3.066000 0.412000 ;
        RECT 2.884000 0.262000 2.945000 0.521000 ;
        RECT 2.811000 0.690000 2.872000 0.888000 ;
        RECT 2.709000 0.152000 2.770000 0.289000 ;
        RECT 2.591000 0.454000 2.652000 0.752000 ;
        RECT 2.516000 0.262000 2.577000 0.399000 ;
        RECT 2.414000 0.807000 2.475000 0.888000 ;
        RECT 2.292000 0.698000 2.353000 1.008000 ;
        RECT 2.170000 0.563000 2.231000 0.899000 ;
        RECT 2.048000 0.563000 2.109000 0.706000 ;
        RECT 2.039000 0.150000 2.100000 0.618000 ;
        RECT 1.902000 0.226000 1.963000 0.899000 ;
        RECT 1.539000 0.368000 1.600000 0.857000 ;
        RECT 1.427000 0.219000 1.488000 0.423000 ;
        RECT 1.417000 0.619000 1.478000 0.988000 ;
        RECT 1.282000 0.329000 1.343000 0.674000 ;
        RECT 0.875000 0.933000 0.936000 1.050000 ;
        RECT 0.753000 0.795000 0.814000 0.936000 ;
        RECT 0.616000 0.154000 0.677000 0.248000 ;
        RECT 0.464000 0.858000 0.525000 1.050000 ;
        RECT 0.390000 0.369000 0.451000 0.755000 ;
        RECT 0.090000 0.319000 0.151000 0.788000 ;
        RECT 3.855000 0.374000 4.058000 0.429000 ;
        RECT 3.573000 0.821000 3.935000 0.876000 ;
        RECT 3.367000 0.931000 4.058000 0.986000 ;
        RECT 3.116000 0.800000 3.634000 0.855000 ;
        RECT 3.005000 0.357000 3.634000 0.412000 ;
        RECT 2.811000 0.690000 3.512000 0.745000 ;
        RECT 2.709000 0.152000 3.066000 0.207000 ;
        RECT 2.591000 0.943000 3.177000 0.998000 ;
        RECT 2.591000 0.576000 3.370000 0.631000 ;
        RECT 2.516000 0.344000 2.945000 0.399000 ;
        RECT 2.414000 0.807000 2.872000 0.862000 ;
        RECT 2.170000 0.563000 2.453000 0.618000 ;
        RECT 2.039000 0.563000 2.109000 0.618000 ;
        RECT 2.030000 0.150000 2.125000 0.205000 ;
        RECT 1.902000 0.844000 2.231000 0.899000 ;
        RECT 1.427000 0.368000 1.808000 0.423000 ;
        RECT 1.315000 0.219000 1.488000 0.274000 ;
        RECT 1.282000 0.619000 1.478000 0.674000 ;
        RECT 0.875000 0.933000 1.678000 0.988000 ;
        RECT 0.753000 0.795000 1.356000 0.850000 ;
        RECT 0.616000 0.193000 1.193000 0.248000 ;
        RECT 0.609000 0.881000 0.814000 0.936000 ;
        RECT 0.487000 0.302000 0.941000 0.357000 ;
        RECT 0.464000 0.995000 0.936000 1.050000 ;
        RECT 0.419000 0.724000 0.692000 0.779000 ;
        RECT 0.390000 0.700000 0.552000 0.755000 ;
        RECT 0.390000 0.369000 0.562000 0.424000 ;
        RECT 0.103000 0.858000 0.525000 0.913000 ;
        RECT 2.884000 0.467000 3.512000 0.521000 ;
        RECT 2.678000 0.235000 2.770000 0.289000 ;
        RECT 2.292000 0.698000 2.681000 0.752000 ;
        RECT 2.161000 0.454000 2.652000 0.508000 ;
        RECT 1.588000 0.954000 2.353000 1.008000 ;
        RECT 0.382000 0.154000 0.677000 0.208000 ;
        RECT 2.048000 0.150000 2.100000 0.706000 ;
        RECT 0.103000 0.319000 0.151000 0.913000 ;
        RECT 0.419000 0.369000 0.451000 0.779000 ;
    END
END SDFFHQX2

MACRO OR4X4
    CLASS CORE ;
    FOREIGN OR4X4 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 2.000000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.683000 0.549000 0.882000 0.639000 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.405000 0.415000 0.592000 0.523000 ;
        RECT 0.937000 0.400000 1.030000 0.494000 ;
        RECT 0.499000 0.415000 0.592000 0.602000 ;
        RECT 0.405000 0.415000 1.030000 0.494000 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.299000 0.633000 0.401000 0.776000 ;
        RECT 0.303000 0.620000 0.397000 0.776000 ;
        RECT 1.128000 0.548000 1.222000 0.629000 ;
        RECT 0.934000 0.700000 1.207000 0.776000 ;
        RECT 0.299000 0.700000 0.423000 0.776000 ;
        RECT 1.143000 0.548000 1.207000 0.776000 ;
        RECT 0.299000 0.721000 1.207000 0.776000 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.220000 0.833000 0.424000 0.926000 ;
        RECT 1.178000 0.388000 1.271000 0.469000 ;
        RECT 0.129000 0.620000 0.193000 0.894000 ;
        RECT 1.302000 0.414000 1.365000 0.888000 ;
        RECT 0.129000 0.833000 0.424000 0.894000 ;
        RECT 1.178000 0.414000 1.365000 0.469000 ;
        RECT 0.129000 0.833000 1.365000 0.888000 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 2.000000 1.280000 ;
        RECT 1.394000 1.078000 1.488000 1.280000 ;
        RECT 1.791000 1.078000 1.884000 1.280000 ;
        RECT 0.050000 0.977000 0.143000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 2.000000 0.080000 ;
        RECT 1.292000 -0.080000 1.386000 0.122000 ;
        RECT 0.457000 -0.080000 0.551000 0.122000 ;
        RECT 1.769000 -0.080000 1.862000 0.122000 ;
        RECT 0.050000 -0.080000 0.143000 0.399000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.493000 0.344000 1.675000 0.793000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.713000 0.154000 0.807000 0.346000 ;
        RECT 0.248000 0.221000 0.342000 0.414000 ;
        RECT 1.758000 0.500000 1.851000 0.581000 ;
        RECT 0.711000 0.944000 0.804000 1.025000 ;
        RECT 1.773000 0.223000 1.836000 0.999000 ;
        RECT 0.566000 0.223000 0.629000 0.345000 ;
        RECT 0.711000 0.944000 1.836000 0.999000 ;
        RECT 0.248000 0.290000 0.629000 0.345000 ;
        RECT 0.566000 0.223000 1.836000 0.277000 ;
    END
END OR4X4

MACRO OR4X2
    CLASS CORE ;
    FOREIGN OR4X2 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.100000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.039000 0.433000 0.151000 0.567000 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.222000 0.167000 0.364000 0.264000 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.406000 0.527000 0.556000 0.633000 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.664000 0.700000 0.878000 0.767000 ;
        RECT 0.664000 0.552000 0.728000 0.767000 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 1.100000 1.280000 ;
        RECT 0.742000 1.078000 0.836000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 1.100000 0.080000 ;
        RECT 0.551000 -0.080000 0.646000 0.122000 ;
        RECT 0.050000 -0.080000 0.144000 0.122000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.942000 0.182000 1.061000 0.375000 ;
        RECT 0.953000 0.700000 1.061000 1.010000 ;
        RECT 0.997000 0.182000 1.061000 1.010000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.812000 0.462000 0.918000 0.576000 ;
        RECT 0.050000 0.731000 0.144000 0.924000 ;
        RECT 0.575000 0.320000 0.669000 0.401000 ;
        RECT 0.215000 0.320000 0.285000 0.388000 ;
        RECT 0.812000 0.333000 0.876000 0.576000 ;
        RECT 0.215000 0.320000 0.279000 0.717000 ;
        RECT 0.081000 0.662000 0.144000 0.924000 ;
        RECT 0.285000 0.333000 0.876000 0.388000 ;
        RECT 0.081000 0.662000 0.279000 0.717000 ;
    END
END OR4X2

MACRO OR4X1
    CLASS CORE ;
    FOREIGN OR4X1 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.100000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.039000 0.656000 0.156000 0.773000 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.222000 0.517000 0.356000 0.635000 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.406000 0.693000 0.550000 0.767000 ;
        RECT 0.486000 0.555000 0.550000 0.767000 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.754000 0.555000 0.886000 0.665000 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 1.100000 1.280000 ;
        RECT 0.689000 1.078000 0.783000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 1.100000 0.080000 ;
        RECT 0.739000 -0.080000 0.833000 0.122000 ;
        RECT 0.217000 -0.080000 0.311000 0.122000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.900000 0.833000 1.061000 0.921000 ;
        RECT 0.950000 0.226000 1.056000 0.307000 ;
        RECT 0.992000 0.226000 1.056000 0.921000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.625000 0.394000 0.915000 0.477000 ;
        RECT 0.572000 0.281000 0.689000 0.362000 ;
        RECT 0.128000 0.343000 0.222000 0.424000 ;
        RECT 0.056000 0.864000 0.150000 0.945000 ;
        RECT 0.625000 0.281000 0.689000 0.932000 ;
        RECT 0.158000 0.281000 0.222000 0.424000 ;
        RECT 0.158000 0.281000 0.689000 0.336000 ;
        RECT 0.056000 0.877000 0.689000 0.932000 ;
    END
END OR4X1

MACRO OR3X4
    CLASS CORE ;
    FOREIGN OR3X4 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.600000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.392000 0.567000 0.548000 0.694000 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.667000 0.457000 0.758000 0.583000 ;
        RECT 0.172000 0.431000 0.264000 0.512000 ;
        RECT 0.172000 0.439000 0.298000 0.512000 ;
        RECT 0.172000 0.457000 0.758000 0.512000 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.038000 0.681000 0.215000 0.775000 ;
        RECT 0.124000 0.604000 0.215000 0.775000 ;
        RECT 0.154000 0.700000 0.236000 0.804000 ;
        RECT 0.038000 0.700000 0.236000 0.775000 ;
        RECT 0.634000 0.704000 0.769000 0.767000 ;
        RECT 0.855000 0.413000 0.917000 0.758000 ;
        RECT 0.634000 0.704000 0.696000 0.804000 ;
        RECT 0.154000 0.604000 0.215000 0.804000 ;
        RECT 0.831000 0.700000 0.917000 0.758000 ;
        RECT 0.855000 0.413000 0.966000 0.468000 ;
        RECT 0.154000 0.749000 0.696000 0.804000 ;
        RECT 0.634000 0.704000 0.917000 0.758000 ;
        END
    END C
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 1.600000 1.280000 ;
        RECT 1.418000 0.983000 1.510000 1.280000 ;
        RECT 1.061000 0.983000 1.153000 1.280000 ;
        RECT 0.048000 1.078000 0.140000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 1.600000 0.080000 ;
        RECT 1.403000 -0.080000 1.495000 0.122000 ;
        RECT 0.529000 -0.080000 0.621000 0.222000 ;
        RECT 0.958000 -0.080000 1.049000 0.122000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.104000 0.331000 1.207000 0.767000 ;
        RECT 1.104000 0.679000 1.339000 0.767000 ;
        RECT 1.104000 0.331000 1.274000 0.412000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.739000 0.213000 0.835000 0.358000 ;
        RECT 0.739000 0.162000 0.831000 0.358000 ;
        RECT 0.322000 0.162000 0.413000 0.358000 ;
        RECT 1.332000 0.532000 1.463000 0.613000 ;
        RECT 0.555000 0.896000 0.646000 0.977000 ;
        RECT 1.401000 0.213000 1.463000 0.898000 ;
        RECT 0.791000 0.843000 0.853000 0.951000 ;
        RECT 0.835000 0.213000 1.463000 0.268000 ;
        RECT 0.791000 0.843000 1.463000 0.898000 ;
        RECT 0.739000 0.213000 1.332000 0.268000 ;
        RECT 0.555000 0.896000 0.853000 0.951000 ;
        RECT 0.322000 0.304000 0.835000 0.358000 ;
    END
END OR3X4

MACRO OR3X1
    CLASS CORE ;
    FOREIGN OR3X1 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.100000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.196000 0.567000 0.336000 0.698000 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.371000 0.412000 0.511000 0.512000 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.544000 0.612000 0.694000 0.767000 ;
        END
    END C
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 1.100000 1.280000 ;
        RECT 0.654000 1.078000 0.749000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 1.100000 0.080000 ;
        RECT 0.286000 -0.080000 0.381000 0.122000 ;
        RECT 0.656000 -0.080000 0.750000 0.122000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.932000 0.555000 1.062000 0.706000 ;
        RECT 0.881000 0.685000 0.996000 0.877000 ;
        RECT 0.903000 0.252000 0.996000 0.337000 ;
        RECT 0.903000 0.252000 0.997000 0.333000 ;
        RECT 0.932000 0.252000 0.996000 0.877000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.046000 0.790000 0.200000 0.877000 ;
        RECT 0.731000 0.286000 0.814000 0.502000 ;
        RECT 0.461000 0.274000 0.556000 0.357000 ;
        RECT 0.046000 0.274000 0.150000 0.357000 ;
        RECT 0.731000 0.421000 0.856000 0.502000 ;
        RECT 0.150000 0.286000 0.814000 0.357000 ;
        RECT 0.046000 0.286000 0.556000 0.357000 ;
        RECT 0.046000 0.274000 0.110000 0.877000 ;
    END
END OR3X1

MACRO OR2X4
    CLASS CORE ;
    FOREIGN OR2X4 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.100000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.039000 0.392000 0.144000 0.556000 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.343000 0.479000 0.511000 0.663000 ;
        END
    END B
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 1.100000 1.280000 ;
        RECT 0.794000 1.078000 0.889000 1.280000 ;
        RECT 0.417000 1.078000 0.511000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 1.100000 0.080000 ;
        RECT 0.461000 -0.080000 0.556000 0.214000 ;
        RECT 0.828000 -0.080000 0.922000 0.122000 ;
        RECT 0.050000 -0.080000 0.144000 0.290000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.589000 0.300000 0.694000 0.633000 ;
        RECT 0.606000 0.624000 0.696000 0.733000 ;
        RECT 0.606000 0.300000 0.694000 0.733000 ;
        RECT 0.606000 0.652000 0.700000 0.733000 ;
        RECT 0.589000 0.324000 0.733000 0.405000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.772000 0.500000 0.867000 0.581000 ;
        RECT 0.214000 0.276000 0.344000 0.357000 ;
        RECT 0.050000 0.669000 0.278000 0.750000 ;
        RECT 0.772000 0.500000 0.836000 0.843000 ;
        RECT 0.214000 0.276000 0.278000 0.843000 ;
        RECT 0.214000 0.788000 0.836000 0.843000 ;
    END
END OR2X4

MACRO OR2X2
    CLASS CORE ;
    FOREIGN OR2X2 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 0.700000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.037000 0.393000 0.138000 0.544000 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.212000 0.414000 0.337000 0.558000 ;
        END
    END B
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 0.700000 1.280000 ;
        RECT 0.345000 1.078000 0.435000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 0.700000 0.080000 ;
        RECT 0.345000 -0.080000 0.435000 0.122000 ;
        RECT 0.048000 -0.080000 0.138000 0.122000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.546000 0.721000 0.650000 0.914000 ;
        RECT 0.548000 0.196000 0.650000 0.389000 ;
        RECT 0.589000 0.196000 0.650000 0.914000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.399000 0.502000 0.528000 0.583000 ;
        RECT 0.196000 0.252000 0.286000 0.333000 ;
        RECT 0.048000 0.721000 0.138000 0.802000 ;
        RECT 0.399000 0.279000 0.460000 0.776000 ;
        RECT 0.048000 0.721000 0.460000 0.776000 ;
        RECT 0.196000 0.279000 0.460000 0.333000 ;
    END
END OR2X2

MACRO OR2X1
    CLASS CORE ;
    FOREIGN OR2X1 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 0.700000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.042000 0.474000 0.154000 0.638000 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.228000 0.567000 0.323000 0.767000 ;
        RECT 0.228000 0.567000 0.313000 0.771000 ;
        RECT 0.212000 0.700000 0.313000 0.771000 ;
        RECT 0.212000 0.700000 0.323000 0.767000 ;
        END
    END B
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 0.700000 1.280000 ;
        RECT 0.290000 1.059000 0.384000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.119000 -0.080000 0.369000 0.122000 ;
        RECT 0.000000 -0.080000 0.700000 0.080000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.562000 0.695000 0.658000 0.867000 ;
        RECT 0.562000 0.314000 0.658000 0.395000 ;
        RECT 0.553000 0.786000 0.658000 0.867000 ;
        RECT 0.597000 0.314000 0.658000 0.867000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.118000 0.313000 0.215000 0.405000 ;
        RECT 0.410000 0.512000 0.536000 0.593000 ;
        RECT 0.053000 0.838000 0.143000 0.919000 ;
        RECT 0.410000 0.313000 0.471000 0.906000 ;
        RECT 0.118000 0.313000 0.471000 0.368000 ;
        RECT 0.053000 0.851000 0.471000 0.906000 ;
    END
END OR2X1

MACRO OAI2BB1X1
    CLASS CORE ;
    FOREIGN OAI2BB1X1 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 0.900000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A0N
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.170000 0.424000 0.322000 0.532000 ;
        END
    END A0N
    PIN A1N
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.038000 0.612000 0.142000 0.767000 ;
        RECT 0.038000 0.612000 0.185000 0.693000 ;
        END
    END A1N
    PIN B0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.398000 0.526000 0.566000 0.640000 ;
        END
    END B0
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.049000 1.078000 0.469000 1.280000 ;
        RECT 0.000000 1.120000 0.900000 1.280000 ;
        RECT 0.738000 1.078000 0.830000 1.280000 ;
        RECT 0.753000 1.065000 0.815000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 0.900000 0.080000 ;
        RECT 0.420000 -0.080000 0.513000 0.122000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.758000 0.343000 0.860000 0.424000 ;
        RECT 0.585000 0.858000 0.678000 0.939000 ;
        RECT 0.779000 0.839000 0.860000 0.913000 ;
        RECT 0.798000 0.343000 0.860000 0.913000 ;
        RECT 0.585000 0.858000 0.860000 0.913000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.213000 0.749000 0.305000 0.843000 ;
        RECT 0.633000 0.500000 0.735000 0.583000 ;
        RECT 0.049000 0.223000 0.142000 0.304000 ;
        RECT 0.633000 0.235000 0.695000 0.804000 ;
        RECT 0.213000 0.749000 0.695000 0.804000 ;
        RECT 0.213000 0.235000 0.695000 0.289000 ;
        RECT 0.142000 0.235000 0.633000 0.289000 ;
        RECT 0.049000 0.235000 0.305000 0.289000 ;
    END
END OAI2BB1X1

MACRO OAI22XL
    CLASS CORE ;
    FOREIGN OAI22XL 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.100000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.575000 0.473000 0.669000 0.652000 ;
        RECT 0.575000 0.573000 0.674000 0.627000 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.772000 0.585000 0.878000 0.767000 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.222000 0.420000 0.444000 0.507000 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.039000 0.639000 0.237000 0.767000 ;
        END
    END B1
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 1.100000 1.280000 ;
        RECT 0.783000 1.078000 0.878000 1.280000 ;
        RECT 0.050000 1.078000 0.144000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 1.100000 0.080000 ;
        RECT 0.261000 -0.080000 0.356000 0.122000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.417000 0.826000 0.511000 0.907000 ;
        RECT 0.672000 0.285000 0.767000 0.365000 ;
        RECT 0.976000 0.387000 1.040000 0.894000 ;
        RECT 0.744000 0.311000 0.808000 0.442000 ;
        RECT 0.744000 0.387000 1.040000 0.442000 ;
        RECT 0.417000 0.839000 1.040000 0.894000 ;
        RECT 0.672000 0.311000 0.808000 0.365000 ;
        RECT 0.744000 0.285000 0.767000 0.442000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.872000 0.251000 0.967000 0.332000 ;
        RECT 0.472000 0.285000 0.567000 0.365000 ;
        RECT 0.872000 0.175000 0.936000 0.332000 ;
        RECT 0.503000 0.175000 0.567000 0.365000 ;
        RECT 0.503000 0.175000 0.936000 0.230000 ;
        RECT 0.050000 0.298000 0.567000 0.352000 ;
    END
END OAI22XL

MACRO OAI22X2
    CLASS CORE ;
    FOREIGN OAI22X2 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.600000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.843000 0.560000 0.948000 0.664000 ;
        RECT 0.843000 0.573000 1.009000 0.664000 ;
        RECT 1.343000 0.583000 1.434000 0.664000 ;
        RECT 0.843000 0.610000 1.434000 0.664000 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.104000 0.412000 1.239000 0.554000 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.048000 0.398000 0.140000 0.554000 ;
        RECT 0.663000 0.473000 0.754000 0.554000 ;
        RECT 0.661000 0.473000 0.754000 0.540000 ;
        RECT 0.661000 0.398000 0.723000 0.540000 ;
        RECT 0.663000 0.398000 0.723000 0.554000 ;
        RECT 0.048000 0.398000 0.723000 0.452000 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.339000 0.508000 0.558000 0.589000 ;
        RECT 0.236000 0.535000 0.298000 0.627000 ;
        RECT 0.236000 0.535000 0.558000 0.589000 ;
        END
    END B1
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 1.600000 1.280000 ;
        RECT 1.096000 0.911000 1.188000 1.280000 ;
        RECT 0.404000 0.911000 0.496000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 1.600000 0.080000 ;
        RECT 0.070000 -0.080000 0.162000 0.122000 ;
        RECT 0.555000 -0.080000 0.646000 0.122000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.441000 0.720000 1.558000 0.833000 ;
        RECT 1.282000 0.746000 1.558000 0.833000 ;
        RECT 1.282000 0.746000 1.364000 0.894000 ;
        RECT 1.309000 0.262000 1.401000 0.343000 ;
        RECT 0.954000 0.262000 1.045000 0.343000 ;
        RECT 0.752000 0.720000 0.843000 0.801000 ;
        RECT 0.048000 0.720000 0.140000 0.801000 ;
        RECT 1.496000 0.288000 1.558000 0.833000 ;
        RECT 0.954000 0.288000 1.558000 0.343000 ;
        RECT 0.048000 0.746000 1.558000 0.801000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.760000 0.261000 0.851000 0.342000 ;
        RECT 0.404000 0.261000 0.496000 0.342000 ;
        RECT 0.048000 0.261000 0.140000 0.342000 ;
        RECT 0.048000 0.287000 0.851000 0.342000 ;
    END
END OAI22X2

MACRO OAI22X1
    CLASS CORE ;
    FOREIGN OAI22X1 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.100000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.575000 0.473000 0.694000 0.633000 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.772000 0.585000 0.878000 0.767000 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.350000 0.433000 0.444000 0.520000 ;
        RECT 0.222000 0.433000 0.444000 0.511000 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.039000 0.567000 0.233000 0.655000 ;
        END
    END B1
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 1.100000 1.280000 ;
        RECT 0.783000 1.078000 0.878000 1.280000 ;
        RECT 0.050000 1.078000 0.144000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 1.100000 0.080000 ;
        RECT 0.261000 -0.080000 0.356000 0.122000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.956000 0.358000 1.040000 0.439000 ;
        RECT 0.672000 0.313000 0.767000 0.394000 ;
        RECT 0.417000 0.826000 0.511000 0.907000 ;
        RECT 0.976000 0.358000 1.040000 0.894000 ;
        RECT 0.703000 0.313000 0.767000 0.413000 ;
        RECT 0.703000 0.358000 1.040000 0.413000 ;
        RECT 0.417000 0.839000 1.040000 0.894000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.872000 0.223000 0.967000 0.304000 ;
        RECT 0.472000 0.298000 0.567000 0.379000 ;
        RECT 0.050000 0.298000 0.144000 0.379000 ;
        RECT 0.872000 0.204000 0.936000 0.304000 ;
        RECT 0.503000 0.204000 0.567000 0.379000 ;
        RECT 0.503000 0.204000 0.936000 0.258000 ;
        RECT 0.144000 0.311000 0.472000 0.365000 ;
    END
END OAI22X1

MACRO OAI221X1
    CLASS CORE ;
    FOREIGN OAI221X1 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.400000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.375000 0.560000 0.581000 0.673000 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.673000 0.567000 0.838000 0.671000 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.212000 0.399000 0.412000 0.500000 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.037000 0.567000 0.223000 0.655000 ;
        END
    END B1
    PIN C0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.017000 0.533000 1.188000 0.640000 ;
        END
    END C0
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 1.400000 1.280000 ;
        RECT 0.748000 1.078000 0.838000 1.280000 ;
        RECT 0.048000 1.078000 0.138000 1.280000 ;
        RECT 0.762000 1.065000 0.823000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 1.400000 0.080000 ;
        RECT 0.451000 -0.080000 0.541000 0.122000 ;
        RECT 0.048000 -0.080000 0.138000 0.122000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.204000 0.282000 1.310000 0.363000 ;
        RECT 0.398000 0.829000 1.358000 0.910000 ;
        RECT 1.249000 0.282000 1.310000 0.910000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 1.013000 0.337000 1.103000 0.418000 ;
        RECT 0.822000 0.226000 0.912000 0.307000 ;
        RECT 0.631000 0.345000 0.721000 0.426000 ;
        RECT 0.249000 0.226000 0.339000 0.307000 ;
        RECT 0.631000 0.363000 1.103000 0.418000 ;
        RECT 0.249000 0.226000 0.912000 0.281000 ;
    END
END OAI221X1

MACRO NOR4BBX2
    CLASS CORE ;
    FOREIGN NOR4BBX2 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 2.000000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN AN
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.160000 0.380000 0.249000 0.500000 ;
        RECT 0.160000 0.433000 0.348000 0.500000 ;
        END
    END AN
    PIN BN
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.556000 0.277000 1.780000 0.396000 ;
        END
    END BN
    PIN C
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.501000 0.457000 0.595000 0.538000 ;
        RECT 0.517000 0.457000 0.595000 0.758000 ;
        RECT 1.315000 0.570000 1.379000 0.758000 ;
        RECT 1.332000 0.704000 1.395000 0.761000 ;
        RECT 1.315000 0.570000 1.416000 0.625000 ;
        RECT 0.517000 0.704000 1.395000 0.758000 ;
        RECT 1.332000 0.570000 1.379000 0.761000 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.315000 0.557000 0.379000 0.876000 ;
        RECT 1.500000 0.570000 1.563000 0.876000 ;
        RECT 0.423000 0.821000 0.486000 0.894000 ;
        RECT 1.500000 0.570000 1.602000 0.625000 ;
        RECT 0.315000 0.821000 1.563000 0.876000 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 2.000000 1.280000 ;
        RECT 0.204000 1.078000 0.298000 1.280000 ;
        RECT 1.590000 1.078000 1.683000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 2.000000 0.080000 ;
        RECT 1.074000 -0.080000 1.168000 0.122000 ;
        RECT 0.248000 -0.080000 0.342000 0.198000 ;
        RECT 0.656000 -0.080000 0.749000 0.122000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.857000 0.894000 1.964000 0.986000 ;
        RECT 0.917000 0.931000 1.032000 1.012000 ;
        RECT 0.865000 0.165000 0.959000 0.246000 ;
        RECT 0.446000 0.165000 0.540000 0.246000 ;
        RECT 1.231000 0.150000 1.295000 0.246000 ;
        RECT 0.968000 0.931000 1.032000 1.027000 ;
        RECT 1.901000 0.150000 1.964000 0.986000 ;
        RECT 1.231000 0.150000 1.964000 0.205000 ;
        RECT 0.917000 0.931000 1.964000 0.986000 ;
        RECT 0.446000 0.192000 1.295000 0.246000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.033000 0.683000 0.143000 0.876000 ;
        RECT 0.033000 0.217000 0.143000 0.324000 ;
        RECT 1.138000 0.457000 1.231000 0.538000 ;
        RECT 0.919000 0.457000 1.012000 0.538000 ;
        RECT 0.697000 0.457000 0.791000 0.538000 ;
        RECT 0.727000 0.457000 0.791000 0.649000 ;
        RECT 0.318000 0.269000 0.382000 0.379000 ;
        RECT 1.774000 0.457000 1.837000 0.764000 ;
        RECT 1.358000 0.262000 1.421000 0.512000 ;
        RECT 1.138000 0.457000 1.201000 0.649000 ;
        RECT 0.919000 0.324000 0.982000 0.538000 ;
        RECT 0.033000 0.217000 0.096000 0.876000 ;
        RECT 1.358000 0.262000 1.493000 0.317000 ;
        RECT 1.138000 0.457000 1.837000 0.512000 ;
        RECT 0.727000 0.594000 1.201000 0.649000 ;
        RECT 0.318000 0.324000 0.982000 0.379000 ;
        RECT 0.143000 0.269000 0.382000 0.324000 ;
    END
END NOR4BBX2

MACRO NOR4XL
    CLASS CORE ;
    FOREIGN NOR4XL 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.100000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.811000 0.494000 0.906000 0.617000 ;
        RECT 0.811000 0.439000 0.878000 0.617000 ;
        RECT 0.793000 0.439000 0.878000 0.494000 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.529000 0.433000 0.646000 0.514000 ;
        RECT 0.529000 0.433000 0.593000 0.761000 ;
        RECT 0.426000 0.700000 0.593000 0.761000 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.222000 0.421000 0.440000 0.526000 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.039000 0.550000 0.158000 0.708000 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 1.100000 1.280000 ;
        RECT 0.050000 1.078000 0.144000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 1.100000 0.080000 ;
        RECT 0.956000 -0.080000 1.050000 0.122000 ;
        RECT 0.517000 -0.080000 0.611000 0.122000 ;
        RECT 0.050000 -0.080000 0.144000 0.122000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.785000 0.698000 0.879000 0.890000 ;
        RECT 0.261000 0.269000 1.040000 0.350000 ;
        RECT 0.976000 0.269000 1.040000 0.761000 ;
        RECT 0.785000 0.706000 1.040000 0.761000 ;
        END
    END Y
END NOR4XL

MACRO NOR4X4
    CLASS CORE ;
    FOREIGN NOR4X4 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 3.000000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.691000 0.573000 0.858000 0.679000 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.864000 0.433000 1.999000 0.538000 ;
        RECT 0.512000 0.392000 0.648000 0.494000 ;
        RECT 1.000000 0.392000 1.091000 0.637000 ;
        RECT 0.512000 0.392000 0.603000 0.538000 ;
        RECT 2.352000 0.457000 2.443000 0.538000 ;
        RECT 1.864000 0.392000 1.925000 0.538000 ;
        RECT 1.864000 0.483000 2.443000 0.538000 ;
        RECT 0.512000 0.392000 1.925000 0.446000 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 2.531000 0.476000 2.622000 0.573000 ;
        RECT 1.178000 0.700000 1.262000 0.789000 ;
        RECT 0.362000 0.706000 0.472000 0.789000 ;
        RECT 1.626000 0.502000 1.754000 0.583000 ;
        RECT 1.201000 0.502000 1.291000 0.583000 ;
        RECT 0.333000 0.556000 0.424000 0.637000 ;
        RECT 0.362000 0.556000 0.424000 0.789000 ;
        RECT 2.531000 0.476000 2.592000 0.648000 ;
        RECT 1.693000 0.502000 1.754000 0.648000 ;
        RECT 1.201000 0.502000 1.262000 0.789000 ;
        RECT 1.693000 0.593000 2.592000 0.648000 ;
        RECT 1.201000 0.502000 1.754000 0.557000 ;
        RECT 0.362000 0.735000 1.262000 0.789000 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.425000 0.618000 1.516000 0.758000 ;
        RECT 2.710000 0.429000 2.809000 0.510000 ;
        RECT 0.055000 0.556000 0.237000 0.637000 ;
        RECT 1.425000 0.618000 1.487000 0.899000 ;
        RECT 0.175000 0.556000 0.237000 0.899000 ;
        RECT 2.710000 0.429000 2.771000 0.758000 ;
        RECT 0.175000 0.844000 1.487000 0.899000 ;
        RECT 1.425000 0.704000 2.771000 0.758000 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 3.000000 1.280000 ;
        RECT 1.432000 1.078000 1.523000 1.280000 ;
        RECT 0.048000 1.078000 0.139000 1.280000 ;
        RECT 2.816000 1.078000 2.906000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 3.000000 0.080000 ;
        RECT 2.424000 -0.080000 2.515000 0.212000 ;
        RECT 2.037000 -0.080000 2.128000 0.212000 ;
        RECT 0.834000 -0.080000 0.925000 0.212000 ;
        RECT 0.440000 -0.080000 0.531000 0.211000 ;
        RECT 0.048000 -0.080000 0.139000 0.211000 ;
        RECT 2.816000 -0.080000 2.906000 0.212000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 2.861000 0.567000 2.963000 0.900000 ;
        RECT 2.861000 0.567000 2.943000 0.923000 ;
        RECT 2.619000 0.256000 2.710000 0.337000 ;
        RECT 2.230000 0.256000 2.321000 0.337000 ;
        RECT 2.108000 0.867000 2.199000 0.948000 ;
        RECT 0.755000 0.954000 0.846000 1.035000 ;
        RECT 0.638000 0.256000 0.729000 0.337000 ;
        RECT 0.245000 0.256000 0.336000 0.337000 ;
        RECT 2.881000 0.282000 2.943000 0.923000 ;
        RECT 2.108000 0.867000 2.170000 1.008000 ;
        RECT 2.108000 0.868000 2.943000 0.923000 ;
        RECT 0.245000 0.282000 2.943000 0.337000 ;
        RECT 0.755000 0.954000 2.170000 1.008000 ;
        END
    END Y
END NOR4X4

MACRO NOR4X2
    CLASS CORE ;
    FOREIGN NOR4X2 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.600000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.710000 0.555000 0.878000 0.636000 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.517000 0.439000 0.607000 0.538000 ;
        RECT 1.007000 0.556000 1.099000 0.637000 ;
        RECT 0.516000 0.457000 0.607000 0.538000 ;
        RECT 1.007000 0.444000 1.069000 0.637000 ;
        RECT 0.517000 0.439000 0.653000 0.499000 ;
        RECT 0.517000 0.444000 1.069000 0.499000 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.365000 0.706000 0.475000 0.789000 ;
        RECT 1.145000 0.396000 1.236000 0.477000 ;
        RECT 0.335000 0.556000 0.427000 0.637000 ;
        RECT 1.174000 0.396000 1.236000 0.789000 ;
        RECT 0.365000 0.556000 0.427000 0.789000 ;
        RECT 0.365000 0.735000 1.236000 0.789000 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.325000 0.556000 1.417000 0.637000 ;
        RECT 0.055000 0.556000 0.238000 0.637000 ;
        RECT 1.325000 0.556000 1.387000 0.899000 ;
        RECT 0.176000 0.556000 0.238000 0.899000 ;
        RECT 0.176000 0.844000 1.387000 0.899000 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 1.600000 1.280000 ;
        RECT 1.442000 1.078000 1.534000 1.280000 ;
        RECT 0.048000 1.078000 0.140000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 1.600000 0.080000 ;
        RECT 0.501000 -0.080000 0.593000 0.122000 ;
        RECT 0.048000 -0.080000 0.140000 0.225000 ;
        RECT 0.927000 -0.080000 1.018000 0.122000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.460000 0.894000 1.542000 1.008000 ;
        RECT 0.761000 0.954000 0.853000 1.035000 ;
        RECT 0.722000 0.261000 0.813000 0.342000 ;
        RECT 0.246000 0.261000 0.338000 0.342000 ;
        RECT 1.480000 0.287000 1.542000 1.008000 ;
        RECT 0.246000 0.287000 1.542000 0.342000 ;
        RECT 0.761000 0.954000 1.542000 1.008000 ;
        END
    END Y
END NOR4X2

MACRO NOR4X1
    CLASS CORE ;
    FOREIGN NOR4X1 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.100000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.811000 0.420000 0.906000 0.560000 ;
        RECT 0.793000 0.439000 0.906000 0.494000 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.529000 0.433000 0.626000 0.514000 ;
        RECT 0.529000 0.433000 0.593000 0.761000 ;
        RECT 0.426000 0.700000 0.593000 0.761000 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.243000 0.421000 0.440000 0.519000 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.062000 0.542000 0.156000 0.700000 ;
        RECT 0.062000 0.542000 0.157000 0.623000 ;
        RECT 0.057000 0.573000 0.156000 0.627000 ;
        RECT 0.057000 0.573000 0.157000 0.623000 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 1.100000 1.280000 ;
        RECT 0.050000 1.078000 0.144000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 1.100000 0.080000 ;
        RECT 0.956000 -0.080000 1.050000 0.122000 ;
        RECT 0.517000 -0.080000 0.611000 0.122000 ;
        RECT 0.050000 -0.080000 0.144000 0.122000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.785000 0.698000 0.879000 0.890000 ;
        RECT 0.261000 0.269000 1.040000 0.350000 ;
        RECT 0.976000 0.269000 1.040000 0.761000 ;
        RECT 0.785000 0.706000 1.040000 0.761000 ;
        END
    END Y
END NOR4X1

MACRO NOR3BX4
    CLASS CORE ;
    FOREIGN NOR3BX4 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 2.000000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN AN
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.180000 0.438000 0.284000 0.519000 ;
        RECT 0.220000 0.306000 0.284000 0.519000 ;
        RECT 0.220000 0.306000 0.304000 0.361000 ;
        END
    END AN
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.565000 0.411000 0.668000 0.513000 ;
        RECT 0.565000 0.411000 0.658000 0.514000 ;
        RECT 1.034000 0.520000 1.128000 0.606000 ;
        RECT 1.032000 0.411000 1.098000 0.500000 ;
        RECT 1.034000 0.411000 1.098000 0.606000 ;
        RECT 1.561000 0.523000 1.624000 0.606000 ;
        RECT 1.034000 0.551000 1.624000 0.606000 ;
        RECT 0.565000 0.411000 1.098000 0.465000 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.231000 0.414000 1.455000 0.495000 ;
        RECT 0.366000 0.536000 0.486000 0.617000 ;
        RECT 1.231000 0.301000 1.295000 0.495000 ;
        RECT 0.423000 0.301000 0.486000 0.627000 ;
        RECT 0.423000 0.301000 1.295000 0.356000 ;
        END
    END C
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 2.000000 1.280000 ;
        RECT 0.264000 0.866000 0.358000 1.280000 ;
        RECT 1.295000 0.911000 1.388000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 2.000000 0.080000 ;
        RECT 1.128000 -0.080000 1.222000 0.122000 ;
        RECT 0.708000 -0.080000 0.802000 0.122000 ;
        RECT 0.300000 -0.080000 0.394000 0.198000 ;
        RECT 1.536000 -0.080000 1.629000 0.198000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.857000 0.433000 1.961000 0.852000 ;
        RECT 1.807000 0.771000 1.961000 0.852000 ;
        RECT 1.337000 0.165000 1.431000 0.246000 ;
        RECT 0.917000 0.165000 1.011000 0.246000 ;
        RECT 0.782000 0.812000 0.876000 0.893000 ;
        RECT 0.499000 0.165000 0.592000 0.246000 ;
        RECT 0.968000 0.771000 1.052000 0.839000 ;
        RECT 0.968000 0.771000 1.032000 0.867000 ;
        RECT 1.857000 0.268000 1.920000 0.852000 ;
        RECT 1.368000 0.165000 1.431000 0.323000 ;
        RECT 1.368000 0.268000 1.920000 0.323000 ;
        RECT 0.968000 0.771000 1.961000 0.826000 ;
        RECT 0.782000 0.812000 1.032000 0.867000 ;
        RECT 0.499000 0.192000 1.431000 0.246000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.780000 0.520000 0.879000 0.756000 ;
        RECT 0.050000 0.701000 0.143000 0.790000 ;
        RECT 0.050000 0.198000 0.157000 0.282000 ;
        RECT 1.687000 0.377000 1.769000 0.715000 ;
        RECT 0.050000 0.198000 0.113000 0.790000 ;
        RECT 1.667000 0.377000 1.769000 0.437000 ;
        RECT 0.050000 0.701000 0.879000 0.756000 ;
        RECT 0.780000 0.661000 1.769000 0.715000 ;
    END
END NOR3BX4

MACRO NOR3BX1
    CLASS CORE ;
    FOREIGN NOR3BX1 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.100000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN AN
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.182000 0.376000 0.286000 0.457000 ;
        RECT 0.222000 0.306000 0.286000 0.457000 ;
        RECT 0.222000 0.306000 0.307000 0.361000 ;
        END
    END AN
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.553000 0.414000 0.756000 0.511000 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.307000 0.536000 0.489000 0.627000 ;
        RECT 0.307000 0.573000 0.490000 0.627000 ;
        END
    END C
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 1.100000 1.280000 ;
        RECT 0.267000 0.897000 0.361000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 1.100000 0.080000 ;
        RECT 0.697000 -0.080000 0.792000 0.122000 ;
        RECT 0.321000 -0.080000 0.415000 0.122000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.783000 0.839000 0.878000 0.924000 ;
        RECT 0.486000 0.269000 1.067000 0.350000 ;
        RECT 1.003000 0.269000 1.067000 0.894000 ;
        RECT 0.783000 0.839000 1.067000 0.894000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.050000 0.237000 0.150000 0.321000 ;
        RECT 0.822000 0.536000 0.917000 0.617000 ;
        RECT 0.050000 0.670000 0.144000 0.751000 ;
        RECT 0.822000 0.536000 0.886000 0.751000 ;
        RECT 0.050000 0.237000 0.114000 0.751000 ;
        RECT 0.050000 0.696000 0.886000 0.751000 ;
    END
END NOR3BX1

MACRO NOR3X4
    CLASS CORE ;
    FOREIGN NOR3X4 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.800000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.638000 0.379000 0.731000 0.496000 ;
        RECT 1.489000 0.581000 1.582000 0.662000 ;
        RECT 0.599000 0.429000 0.731000 0.494000 ;
        RECT 1.490000 0.379000 1.553000 0.662000 ;
        RECT 0.638000 0.379000 1.553000 0.433000 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.311000 0.507000 0.404000 0.610000 ;
        RECT 0.908000 0.488000 0.971000 0.610000 ;
        RECT 0.311000 0.439000 0.374000 0.610000 ;
        RECT 0.908000 0.488000 1.390000 0.543000 ;
        RECT 0.311000 0.555000 0.971000 0.610000 ;
        RECT 0.239000 0.439000 0.374000 0.494000 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.092000 0.598000 1.189000 0.774000 ;
        RECT 0.056000 0.526000 0.153000 0.627000 ;
        RECT 1.021000 0.700000 1.189000 0.774000 ;
        RECT 0.090000 0.526000 0.153000 0.774000 ;
        RECT 0.090000 0.719000 1.189000 0.774000 ;
        END
    END C
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 1.800000 1.280000 ;
        RECT 1.088000 0.989000 1.181000 1.280000 ;
        RECT 0.049000 0.929000 0.142000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 1.800000 0.080000 ;
        RECT 1.227000 -0.080000 1.320000 0.198000 ;
        RECT 0.442000 -0.080000 0.535000 0.198000 ;
        RECT 0.049000 -0.080000 0.142000 0.211000 ;
        RECT 0.835000 -0.080000 0.927000 0.198000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.658000 0.567000 1.762000 0.900000 ;
        RECT 1.561000 0.810000 1.762000 0.892000 ;
        RECT 1.031000 0.242000 1.124000 0.323000 ;
        RECT 0.638000 0.242000 0.731000 0.323000 ;
        RECT 0.573000 0.837000 0.665000 0.918000 ;
        RECT 0.245000 0.242000 0.338000 0.323000 ;
        RECT 1.658000 0.268000 1.721000 0.900000 ;
        RECT 0.573000 0.837000 1.762000 0.892000 ;
        RECT 0.245000 0.268000 1.721000 0.323000 ;
        END
    END Y
END NOR3X4

MACRO NOR3X2
    CLASS CORE ;
    FOREIGN NOR3X2 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.300000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.498000 0.439000 0.682000 0.525000 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.321000 0.445000 0.415000 0.539000 ;
        RECT 0.847000 0.377000 0.943000 0.458000 ;
        RECT 0.321000 0.458000 0.416000 0.539000 ;
        RECT 0.848000 0.377000 0.913000 0.635000 ;
        RECT 0.352000 0.458000 0.416000 0.635000 ;
        RECT 0.352000 0.445000 0.415000 0.635000 ;
        RECT 0.246000 0.439000 0.311000 0.500000 ;
        RECT 0.352000 0.580000 0.913000 0.635000 ;
        RECT 0.246000 0.445000 0.415000 0.500000 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.118000 0.573000 0.214000 0.707000 ;
        RECT 1.007000 0.537000 1.088000 0.744000 ;
        RECT 0.149000 0.573000 0.214000 0.744000 ;
        RECT 0.149000 0.689000 1.088000 0.744000 ;
        RECT 0.058000 0.573000 0.214000 0.627000 ;
        END
    END C
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 1.300000 1.280000 ;
        RECT 1.109000 0.925000 1.204000 1.280000 ;
        RECT 0.051000 0.876000 0.146000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 1.300000 0.080000 ;
        RECT 0.456000 -0.080000 0.552000 0.211000 ;
        RECT 0.051000 -0.080000 0.146000 0.211000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.658000 0.151000 0.754000 0.344000 ;
        RECT 0.253000 0.151000 0.349000 0.344000 ;
        RECT 0.591000 0.800000 0.687000 0.890000 ;
        RECT 1.154000 0.767000 1.240000 0.855000 ;
        RECT 1.175000 0.255000 1.240000 0.855000 ;
        RECT 0.658000 0.255000 1.240000 0.310000 ;
        RECT 0.591000 0.800000 1.240000 0.855000 ;
        RECT 0.253000 0.289000 0.754000 0.344000 ;
        END
    END Y
END NOR3X2

MACRO NOR3X1
    CLASS CORE ;
    FOREIGN NOR3X1 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 0.700000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.456000 0.536000 0.546000 0.617000 ;
        RECT 0.456000 0.536000 0.517000 0.761000 ;
        RECT 0.407000 0.706000 0.517000 0.761000 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.232000 0.421000 0.361000 0.561000 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.048000 0.536000 0.137000 0.694000 ;
        RECT 0.048000 0.536000 0.138000 0.617000 ;
        END
    END C
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 0.700000 1.280000 ;
        RECT 0.048000 0.900000 0.138000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 0.700000 0.080000 ;
        RECT 0.345000 -0.080000 0.435000 0.122000 ;
        RECT 0.048000 -0.080000 0.138000 0.122000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.557000 0.839000 0.666000 0.924000 ;
        RECT 0.196000 0.269000 0.668000 0.350000 ;
        RECT 0.607000 0.269000 0.668000 0.894000 ;
        RECT 0.607000 0.269000 0.666000 0.924000 ;
        RECT 0.557000 0.839000 0.668000 0.894000 ;
        END
    END Y
END NOR3X1

MACRO NOR2BX4
    CLASS CORE ;
    FOREIGN NOR2BX4 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.400000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN AN
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.034000 0.436000 0.138000 0.571000 ;
        END
    END AN
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.321000 0.521000 0.411000 0.650000 ;
        RECT 0.936000 0.563000 1.026000 0.650000 ;
        RECT 0.321000 0.565000 0.468000 0.650000 ;
        RECT 0.321000 0.595000 1.026000 0.650000 ;
        END
    END B
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.223000 1.117000 1.013000 1.280000 ;
        RECT 0.000000 1.120000 1.400000 1.280000 ;
        RECT 0.923000 1.078000 1.013000 1.280000 ;
        RECT 0.223000 1.078000 0.313000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 1.400000 0.080000 ;
        RECT 0.681000 -0.080000 0.772000 0.122000 ;
        RECT 1.087000 -0.080000 1.177000 0.122000 ;
        RECT 0.276000 -0.080000 0.366000 0.122000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.262000 0.264000 1.363000 0.786000 ;
        RECT 1.252000 0.693000 1.363000 0.786000 ;
        RECT 0.883000 0.255000 0.973000 0.336000 ;
        RECT 0.573000 0.705000 1.363000 0.786000 ;
        RECT 0.480000 0.255000 0.570000 0.336000 ;
        RECT 0.883000 0.264000 1.363000 0.336000 ;
        RECT 0.480000 0.281000 1.363000 0.336000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.578000 0.392000 0.668000 0.538000 ;
        RECT 0.074000 0.281000 0.164000 0.362000 ;
        RECT 0.048000 0.793000 0.138000 0.874000 ;
        RECT 1.139000 0.392000 1.200000 0.546000 ;
        RECT 0.199000 0.307000 0.260000 0.848000 ;
        RECT 0.074000 0.307000 0.260000 0.362000 ;
        RECT 0.048000 0.793000 0.260000 0.848000 ;
        RECT 0.578000 0.392000 1.200000 0.446000 ;
        RECT 0.260000 0.392000 0.578000 0.446000 ;
    END
END NOR2BX4

MACRO NOR2BX1
    CLASS CORE ;
    FOREIGN NOR2BX1 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 0.700000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN AN
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.037000 0.486000 0.138000 0.633000 ;
        END
    END AN
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.321000 0.567000 0.411000 0.670000 ;
        RECT 0.321000 0.567000 0.525000 0.633000 ;
        END
    END B
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 0.700000 1.280000 ;
        RECT 0.212000 0.916000 0.302000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 0.700000 0.080000 ;
        RECT 0.562000 -0.080000 0.652000 0.122000 ;
        RECT 0.263000 -0.080000 0.353000 0.122000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.562000 0.706000 0.666000 0.858000 ;
        RECT 0.411000 0.269000 0.501000 0.350000 ;
        RECT 0.605000 0.295000 0.666000 0.858000 ;
        RECT 0.411000 0.295000 0.666000 0.350000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.461000 0.430000 0.544000 0.511000 ;
        RECT 0.048000 0.715000 0.138000 0.796000 ;
        RECT 0.048000 0.304000 0.138000 0.385000 ;
        RECT 0.048000 0.323000 0.260000 0.385000 ;
        RECT 0.199000 0.323000 0.260000 0.770000 ;
        RECT 0.260000 0.443000 0.461000 0.498000 ;
        RECT 0.048000 0.715000 0.260000 0.770000 ;
    END
END NOR2BX1

MACRO NOR2XL
    CLASS CORE ;
    FOREIGN NOR2XL 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 0.600000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.242000 0.406000 0.421000 0.502000 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.061000 0.548000 0.164000 0.633000 ;
        RECT 0.042000 0.567000 0.255000 0.633000 ;
        END
    END B
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 0.600000 1.280000 ;
        RECT 0.055000 1.078000 0.158000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 0.600000 0.080000 ;
        RECT 0.442000 -0.080000 0.545000 0.122000 ;
        RECT 0.055000 -0.080000 0.158000 0.122000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.442000 0.626000 0.561000 0.774000 ;
        RECT 0.248000 0.269000 0.352000 0.350000 ;
        RECT 0.491000 0.295000 0.561000 0.774000 ;
        RECT 0.248000 0.295000 0.561000 0.350000 ;
        END
    END Y
END NOR2XL

MACRO NOR2X4
    CLASS CORE ;
    FOREIGN NOR2X4 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.300000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.432000 0.439000 0.523000 0.525000 ;
        RECT 0.990000 0.464000 1.086000 0.545000 ;
        RECT 0.990000 0.394000 1.055000 0.545000 ;
        RECT 0.459000 0.394000 0.523000 0.525000 ;
        RECT 0.459000 0.394000 1.055000 0.449000 ;
        RECT 0.428000 0.470000 0.523000 0.525000 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.763000 0.561000 0.858000 0.642000 ;
        RECT 0.138000 0.492000 0.234000 0.573000 ;
        RECT 0.246000 0.650000 0.311000 0.761000 ;
        RECT 0.169000 0.492000 0.234000 0.707000 ;
        RECT 0.763000 0.561000 0.827000 0.705000 ;
        RECT 0.169000 0.650000 0.311000 0.707000 ;
        RECT 0.169000 0.650000 0.827000 0.705000 ;
        END
    END B
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 1.300000 1.280000 ;
        RECT 0.799000 1.078000 0.895000 1.280000 ;
        RECT 0.056000 1.078000 0.152000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 1.300000 0.080000 ;
        RECT 0.467000 -0.080000 0.563000 0.211000 ;
        RECT 0.884000 -0.080000 0.979000 0.122000 ;
        RECT 0.051000 -0.080000 0.146000 0.298000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.154000 0.433000 1.261000 0.767000 ;
        RECT 1.148000 0.693000 1.244000 0.840000 ;
        RECT 1.154000 0.433000 1.244000 0.840000 ;
        RECT 1.165000 0.265000 1.249000 0.767000 ;
        RECT 0.670000 0.256000 0.765000 0.337000 ;
        RECT 0.265000 0.256000 0.360000 0.337000 ;
        RECT 0.428000 0.760000 1.244000 0.840000 ;
        RECT 1.165000 0.265000 1.244000 0.840000 ;
        RECT 1.148000 0.693000 1.261000 0.767000 ;
        RECT 0.670000 0.265000 1.249000 0.337000 ;
        RECT 0.265000 0.282000 1.249000 0.337000 ;
        END
    END Y
END NOR2X4

MACRO NOR2X2
    CLASS CORE ;
    FOREIGN NOR2X2 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 0.900000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.327000 0.538000 0.502000 0.633000 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.120000 0.418000 0.229000 0.518000 ;
        RECT 0.652000 0.418000 0.742000 0.564000 ;
        RECT 0.059000 0.418000 0.229000 0.494000 ;
        RECT 0.059000 0.418000 0.742000 0.473000 ;
        END
    END B
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 0.900000 1.280000 ;
        RECT 0.758000 1.078000 0.851000 1.280000 ;
        RECT 0.049000 1.078000 0.142000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 0.900000 0.080000 ;
        RECT 0.758000 -0.080000 0.851000 0.228000 ;
        RECT 0.365000 -0.080000 0.458000 0.340000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.562000 0.170000 0.655000 0.363000 ;
        RECT 0.404000 0.712000 0.496000 0.793000 ;
        RECT 0.805000 0.308000 0.867000 0.761000 ;
        RECT 0.779000 0.706000 0.862000 0.767000 ;
        RECT 0.805000 0.308000 0.862000 0.767000 ;
        RECT 0.779000 0.706000 0.867000 0.761000 ;
        RECT 0.562000 0.308000 0.867000 0.363000 ;
        RECT 0.404000 0.712000 0.862000 0.767000 ;
        END
    END Y
END NOR2X2

MACRO NOR2X1
    CLASS CORE ;
    FOREIGN NOR2X1 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 0.600000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.242000 0.407000 0.421000 0.502000 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.061000 0.548000 0.164000 0.643000 ;
        RECT 0.042000 0.567000 0.255000 0.643000 ;
        END
    END B
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 0.600000 1.280000 ;
        RECT 0.055000 1.078000 0.158000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 0.600000 0.080000 ;
        RECT 0.442000 -0.080000 0.545000 0.122000 ;
        RECT 0.055000 -0.080000 0.158000 0.122000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.442000 0.626000 0.561000 0.774000 ;
        RECT 0.248000 0.269000 0.352000 0.350000 ;
        RECT 0.491000 0.295000 0.561000 0.774000 ;
        RECT 0.248000 0.295000 0.561000 0.350000 ;
        END
    END Y
END NOR2X1

MACRO NAND4BX4
    CLASS CORE ;
    FOREIGN NAND4BX4 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 3.200000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN AN
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.042000 0.433000 0.144000 0.574000 ;
        END
    END AN
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 2.349000 0.433000 2.451000 0.596000 ;
        RECT 2.003000 0.510000 2.104000 0.596000 ;
        RECT 1.121000 0.510000 1.222000 0.596000 ;
        RECT 2.349000 0.515000 2.465000 0.596000 ;
        RECT 0.723000 0.515000 0.824000 0.596000 ;
        RECT 2.003000 0.542000 2.465000 0.596000 ;
        RECT 1.121000 0.510000 2.104000 0.564000 ;
        RECT 0.723000 0.542000 1.222000 0.596000 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 2.591000 0.519000 2.683000 0.600000 ;
        RECT 1.825000 0.625000 1.916000 0.706000 ;
        RECT 1.309000 0.625000 1.401000 0.706000 ;
        RECT 0.544000 0.519000 0.653000 0.600000 ;
        RECT 2.591000 0.519000 2.668000 0.633000 ;
        RECT 2.527000 0.579000 2.589000 0.706000 ;
        RECT 0.591000 0.519000 0.653000 0.706000 ;
        RECT 2.547000 0.573000 2.668000 0.633000 ;
        RECT 1.825000 0.651000 2.589000 0.706000 ;
        RECT 1.309000 0.625000 1.916000 0.680000 ;
        RECT 0.591000 0.651000 1.401000 0.706000 ;
        RECT 2.527000 0.579000 2.668000 0.633000 ;
        RECT 2.547000 0.573000 2.589000 0.706000 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 2.769000 0.426000 2.859000 0.507000 ;
        RECT 0.361000 0.519000 0.453000 0.600000 ;
        RECT 1.568000 0.735000 1.659000 0.815000 ;
        RECT 2.753000 0.439000 2.859000 0.507000 ;
        RECT 2.753000 0.439000 2.815000 0.815000 ;
        RECT 0.413000 0.706000 0.475000 0.815000 ;
        RECT 0.391000 0.519000 0.453000 0.761000 ;
        RECT 0.391000 0.706000 0.475000 0.761000 ;
        RECT 0.413000 0.761000 2.815000 0.815000 ;
        RECT 2.769000 0.426000 2.815000 0.815000 ;
        RECT 0.413000 0.519000 0.453000 0.815000 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 3.200000 1.280000 ;
        RECT 2.078000 1.078000 2.199000 1.280000 ;
        RECT 1.028000 1.078000 1.149000 1.280000 ;
        RECT 2.859000 1.078000 2.951000 1.280000 ;
        RECT 0.276000 1.078000 0.368000 1.280000 ;
        RECT 2.477000 1.078000 2.568000 1.280000 ;
        RECT 0.659000 1.078000 0.750000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 3.200000 0.080000 ;
        RECT 2.882000 -0.080000 2.974000 0.122000 ;
        RECT 0.253000 -0.080000 0.345000 0.122000 ;
        RECT 1.568000 -0.080000 1.659000 0.122000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 2.882000 0.567000 2.985000 0.900000 ;
        RECT 2.882000 0.567000 2.974000 0.942000 ;
        RECT 0.910000 0.150000 1.002000 0.343000 ;
        RECT 2.225000 0.150000 2.316000 0.343000 ;
        RECT 2.294000 0.870000 2.974000 0.942000 ;
        RECT 0.910000 0.207000 2.316000 0.274000 ;
        RECT 0.467000 0.870000 2.974000 0.937000 ;
        RECT 2.921000 0.288000 2.983000 0.900000 ;
        RECT 2.225000 0.288000 2.983000 0.343000 ;
        RECT 2.921000 0.288000 2.974000 0.942000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 2.180000 0.400000 2.281000 0.487000 ;
        RECT 0.909000 0.400000 1.010000 0.487000 ;
        RECT 0.048000 0.801000 0.140000 0.882000 ;
        RECT 0.048000 0.276000 0.140000 0.357000 ;
        RECT 0.210000 0.302000 0.272000 0.856000 ;
        RECT 0.909000 0.400000 2.281000 0.455000 ;
        RECT 0.272000 0.400000 0.909000 0.455000 ;
        RECT 0.048000 0.801000 0.272000 0.856000 ;
        RECT 0.048000 0.302000 0.272000 0.357000 ;
    END
END NAND4BX4

MACRO NAND4BX2
    CLASS CORE ;
    FOREIGN NAND4BX2 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.800000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN AN
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.042000 0.433000 0.146000 0.574000 ;
        END
    END AN
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.085000 0.514000 1.188000 0.596000 ;
        RECT 0.698000 0.515000 0.800000 0.596000 ;
        RECT 1.118000 0.433000 1.188000 0.596000 ;
        RECT 1.118000 0.439000 1.201000 0.494000 ;
        RECT 0.698000 0.542000 1.188000 0.596000 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.285000 0.519000 1.377000 0.627000 ;
        RECT 0.521000 0.519000 0.627000 0.600000 ;
        RECT 1.285000 0.519000 1.347000 0.706000 ;
        RECT 0.565000 0.519000 0.627000 0.706000 ;
        RECT 0.565000 0.651000 1.347000 0.706000 ;
        RECT 1.285000 0.573000 1.381000 0.627000 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.357000 0.761000 1.450000 0.842000 ;
        RECT 0.340000 0.519000 0.424000 0.600000 ;
        RECT 0.361000 0.519000 0.424000 0.761000 ;
        RECT 0.419000 0.706000 0.481000 0.815000 ;
        RECT 0.361000 0.706000 0.481000 0.761000 ;
        RECT 0.419000 0.761000 1.450000 0.815000 ;
        RECT 0.419000 0.519000 0.424000 0.815000 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 1.800000 1.280000 ;
        RECT 1.006000 1.078000 1.129000 1.280000 ;
        RECT 0.245000 1.078000 0.338000 1.280000 ;
        RECT 0.633000 1.078000 0.725000 1.280000 ;
        RECT 0.260000 1.065000 0.323000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 1.800000 0.080000 ;
        RECT 1.560000 -0.080000 1.653000 0.122000 ;
        RECT 0.229000 -0.080000 0.322000 0.122000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.895000 0.150000 0.987000 0.343000 ;
        RECT 1.658000 0.195000 1.741000 0.306000 ;
        RECT 1.658000 0.564000 1.740000 0.973000 ;
        RECT 0.963000 0.870000 1.045000 0.973000 ;
        RECT 1.665000 0.195000 1.741000 0.633000 ;
        RECT 1.665000 0.195000 1.740000 0.973000 ;
        RECT 0.963000 0.901000 1.740000 0.973000 ;
        RECT 0.439000 0.870000 1.045000 0.942000 ;
        RECT 1.658000 0.564000 1.741000 0.633000 ;
        RECT 0.895000 0.195000 1.741000 0.262000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.886000 0.400000 0.989000 0.487000 ;
        RECT 0.049000 0.731000 0.142000 0.812000 ;
        RECT 0.049000 0.276000 0.142000 0.357000 ;
        RECT 0.211000 0.302000 0.274000 0.799000 ;
        RECT 0.274000 0.400000 0.886000 0.455000 ;
        RECT 0.049000 0.744000 0.274000 0.799000 ;
        RECT 0.049000 0.302000 0.274000 0.357000 ;
    END
END NAND4BX2

MACRO NAND4BX1
    CLASS CORE ;
    FOREIGN NAND4BX1 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.300000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN AN
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.950000 0.498000 1.075000 0.633000 ;
        RECT 0.950000 0.498000 1.089000 0.579000 ;
        END
    END AN
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.567000 0.555000 0.743000 0.665000 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.348000 0.555000 0.443000 0.636000 ;
        RECT 0.348000 0.555000 0.466000 0.623000 ;
        RECT 0.401000 0.439000 0.466000 0.623000 ;
        RECT 0.401000 0.439000 0.497000 0.494000 ;
        RECT 0.401000 0.439000 0.443000 0.636000 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.162000 0.492000 0.252000 0.600000 ;
        RECT 0.187000 0.439000 0.252000 0.600000 ;
        RECT 0.187000 0.439000 0.311000 0.494000 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 1.300000 1.280000 ;
        RECT 0.830000 1.078000 0.957000 1.280000 ;
        RECT 0.459000 1.078000 0.554000 1.280000 ;
        RECT 0.079000 1.078000 0.174000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 1.300000 0.080000 ;
        RECT 0.055000 -0.080000 0.151000 0.122000 ;
        RECT 1.154000 -0.080000 1.249000 0.122000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.650000 0.737000 0.746000 0.839000 ;
        RECT 1.154000 0.201000 1.240000 0.306000 ;
        RECT 0.741000 0.201000 0.837000 0.282000 ;
        RECT 0.267000 0.737000 0.363000 0.818000 ;
        RECT 0.597000 0.763000 0.746000 0.839000 ;
        RECT 1.200000 0.573000 1.265000 0.933000 ;
        RECT 1.175000 0.201000 1.240000 0.627000 ;
        RECT 0.681000 0.737000 0.746000 0.933000 ;
        RECT 0.741000 0.201000 1.240000 0.256000 ;
        RECT 0.267000 0.763000 0.746000 0.818000 ;
        RECT 1.175000 0.573000 1.265000 0.627000 ;
        RECT 0.681000 0.879000 1.265000 0.933000 ;
        RECT 1.200000 0.201000 1.240000 0.933000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 1.040000 0.737000 1.135000 0.818000 ;
        RECT 0.938000 0.311000 1.034000 0.392000 ;
        RECT 0.758000 0.419000 0.881000 0.500000 ;
        RECT 0.927000 0.324000 1.034000 0.392000 ;
        RECT 0.927000 0.324000 0.992000 0.405000 ;
        RECT 0.816000 0.350000 0.881000 0.792000 ;
        RECT 0.816000 0.737000 1.135000 0.792000 ;
        RECT 0.816000 0.350000 0.992000 0.405000 ;
        RECT 0.938000 0.311000 0.992000 0.405000 ;
    END
END NAND4BX1

MACRO NAND4X4
    CLASS CORE ;
    FOREIGN NAND4X4 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 3.000000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.988000 0.400000 2.088000 0.487000 ;
        RECT 0.726000 0.400000 0.826000 0.487000 ;
        RECT 0.430000 0.306000 0.492000 0.455000 ;
        RECT 0.430000 0.400000 2.088000 0.455000 ;
        RECT 0.410000 0.306000 0.492000 0.361000 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 2.155000 0.433000 2.257000 0.596000 ;
        RECT 1.811000 0.510000 1.912000 0.596000 ;
        RECT 0.936000 0.510000 1.036000 0.596000 ;
        RECT 2.155000 0.515000 2.270000 0.596000 ;
        RECT 0.541000 0.515000 0.642000 0.596000 ;
        RECT 1.811000 0.542000 2.270000 0.596000 ;
        RECT 0.936000 0.510000 1.912000 0.564000 ;
        RECT 0.541000 0.542000 1.036000 0.596000 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 2.396000 0.519000 2.487000 0.600000 ;
        RECT 1.635000 0.625000 1.726000 0.706000 ;
        RECT 1.123000 0.625000 1.214000 0.706000 ;
        RECT 0.364000 0.519000 0.472000 0.600000 ;
        RECT 2.396000 0.519000 2.472000 0.633000 ;
        RECT 0.410000 0.519000 0.472000 0.706000 ;
        RECT 2.332000 0.579000 2.393000 0.706000 ;
        RECT 2.352000 0.573000 2.472000 0.633000 ;
        RECT 1.635000 0.651000 2.393000 0.706000 ;
        RECT 1.123000 0.625000 1.726000 0.680000 ;
        RECT 0.410000 0.651000 1.214000 0.706000 ;
        RECT 2.332000 0.579000 2.472000 0.633000 ;
        RECT 2.352000 0.573000 2.393000 0.706000 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 2.572000 0.426000 2.662000 0.507000 ;
        RECT 0.182000 0.519000 0.273000 0.600000 ;
        RECT 1.380000 0.735000 1.471000 0.815000 ;
        RECT 2.556000 0.439000 2.662000 0.507000 ;
        RECT 2.556000 0.439000 2.618000 0.815000 ;
        RECT 0.211000 0.519000 0.273000 0.761000 ;
        RECT 0.234000 0.706000 0.295000 0.815000 ;
        RECT 0.211000 0.706000 0.295000 0.761000 ;
        RECT 0.234000 0.761000 2.618000 0.815000 ;
        RECT 2.572000 0.426000 2.618000 0.815000 ;
        RECT 0.234000 0.519000 0.273000 0.815000 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 3.000000 1.280000 ;
        RECT 1.886000 1.078000 2.007000 1.280000 ;
        RECT 0.844000 1.078000 0.964000 1.280000 ;
        RECT 2.662000 1.078000 2.753000 1.280000 ;
        RECT 2.282000 1.078000 2.373000 1.280000 ;
        RECT 0.477000 1.078000 0.568000 1.280000 ;
        RECT 0.098000 1.078000 0.189000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 3.000000 0.080000 ;
        RECT 2.684000 -0.080000 2.775000 0.122000 ;
        RECT 1.380000 -0.080000 1.471000 0.122000 ;
        RECT 0.075000 -0.080000 0.166000 0.122000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 2.684000 0.192000 2.803000 0.307000 ;
        RECT 2.032000 0.150000 2.176000 0.263000 ;
        RECT 2.684000 0.567000 2.786000 0.900000 ;
        RECT 2.684000 0.567000 2.775000 0.942000 ;
        RECT 2.032000 0.150000 2.123000 0.343000 ;
        RECT 0.727000 0.150000 0.818000 0.343000 ;
        RECT 2.723000 0.192000 2.803000 0.639000 ;
        RECT 2.684000 0.567000 2.803000 0.639000 ;
        RECT 2.100000 0.870000 2.775000 0.942000 ;
        RECT 2.032000 0.192000 2.803000 0.263000 ;
        RECT 0.727000 0.207000 2.123000 0.274000 ;
        RECT 0.287000 0.870000 2.775000 0.937000 ;
        RECT 2.723000 0.192000 2.786000 0.900000 ;
        RECT 0.727000 0.207000 2.803000 0.263000 ;
        RECT 2.723000 0.192000 2.775000 0.942000 ;
        END
    END Y
END NAND4X4

MACRO NAND4X2
    CLASS CORE ;
    FOREIGN NAND4X2 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.600000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.698000 0.401000 0.799000 0.487000 ;
        RECT 0.434000 0.306000 0.496000 0.456000 ;
        RECT 0.434000 0.401000 0.799000 0.456000 ;
        RECT 0.413000 0.306000 0.496000 0.361000 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.916000 0.439000 1.017000 0.596000 ;
        RECT 0.512000 0.515000 0.613000 0.596000 ;
        RECT 0.512000 0.542000 1.017000 0.596000 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.102000 0.519000 1.187000 0.627000 ;
        RECT 1.102000 0.519000 1.193000 0.600000 ;
        RECT 0.333000 0.519000 0.442000 0.600000 ;
        RECT 1.102000 0.519000 1.164000 0.706000 ;
        RECT 0.380000 0.519000 0.442000 0.706000 ;
        RECT 0.380000 0.651000 1.164000 0.706000 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.162000 0.761000 1.254000 0.842000 ;
        RECT 0.149000 0.519000 0.241000 0.600000 ;
        RECT 0.236000 0.706000 0.298000 0.815000 ;
        RECT 0.179000 0.519000 0.241000 0.761000 ;
        RECT 0.179000 0.706000 0.298000 0.761000 ;
        RECT 0.236000 0.761000 1.254000 0.815000 ;
        RECT 0.236000 0.519000 0.241000 0.815000 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 1.600000 1.280000 ;
        RECT 0.816000 1.078000 0.937000 1.280000 ;
        RECT 0.447000 1.078000 0.539000 1.280000 ;
        RECT 0.065000 1.078000 0.156000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 1.600000 0.080000 ;
        RECT 1.363000 -0.080000 1.455000 0.122000 ;
        RECT 0.048000 -0.080000 0.140000 0.122000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.706000 0.150000 0.797000 0.343000 ;
        RECT 1.460000 0.195000 1.542000 0.306000 ;
        RECT 1.460000 0.564000 1.541000 0.973000 ;
        RECT 0.773000 0.870000 0.854000 0.973000 ;
        RECT 1.467000 0.195000 1.542000 0.633000 ;
        RECT 1.467000 0.195000 1.541000 0.973000 ;
        RECT 0.773000 0.901000 1.541000 0.973000 ;
        RECT 0.256000 0.870000 0.854000 0.942000 ;
        RECT 1.460000 0.564000 1.542000 0.633000 ;
        RECT 0.706000 0.195000 1.542000 0.262000 ;
        END
    END Y
END NAND4X2

MACRO NAND4X1
    CLASS CORE ;
    FOREIGN NAND4X1 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 0.900000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.645000 0.419000 0.738000 0.500000 ;
        RECT 0.419000 0.439000 0.738000 0.494000 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.521000 0.573000 0.682000 0.662000 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.273000 0.555000 0.405000 0.636000 ;
        RECT 0.273000 0.439000 0.335000 0.636000 ;
        RECT 0.239000 0.439000 0.335000 0.494000 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.079000 0.555000 0.210000 0.636000 ;
        RECT 0.079000 0.439000 0.142000 0.636000 ;
        RECT 0.059000 0.439000 0.142000 0.494000 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 0.900000 1.280000 ;
        RECT 0.758000 1.078000 0.851000 1.280000 ;
        RECT 0.049000 1.078000 0.142000 1.280000 ;
        RECT 0.475000 1.078000 0.567000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 0.900000 0.080000 ;
        RECT 0.053000 -0.080000 0.146000 0.247000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.724000 0.170000 0.817000 0.363000 ;
        RECT 0.758000 0.706000 0.865000 0.792000 ;
        RECT 0.589000 0.737000 0.682000 0.818000 ;
        RECT 0.218000 0.737000 0.311000 0.818000 ;
        RECT 0.802000 0.308000 0.865000 0.792000 ;
        RECT 0.724000 0.308000 0.865000 0.363000 ;
        RECT 0.218000 0.737000 0.865000 0.792000 ;
        RECT 0.802000 0.170000 0.817000 0.792000 ;
        END
    END Y
END NAND4X1

MACRO NAND3BX2
    CLASS CORE ;
    FOREIGN NAND3BX2 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.400000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN AN
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.262000 0.467000 1.363000 0.594000 ;
        RECT 1.267000 0.433000 1.358000 0.594000 ;
        END
    END AN
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.737000 0.433000 0.838000 0.604000 ;
        RECT 0.355000 0.514000 0.445000 0.604000 ;
        RECT 0.737000 0.507000 0.870000 0.588000 ;
        RECT 0.355000 0.549000 0.838000 0.604000 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.082000 0.439000 0.172000 0.573000 ;
        RECT 0.957000 0.462000 1.047000 0.543000 ;
        RECT 0.972000 0.462000 1.033000 0.881000 ;
        RECT 0.111000 0.439000 0.172000 0.881000 ;
        RECT 0.111000 0.826000 1.033000 0.881000 ;
        RECT 0.057000 0.439000 0.172000 0.494000 ;
        END
    END C
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 1.400000 1.280000 ;
        RECT 1.058000 0.952000 1.148000 1.280000 ;
        RECT 0.471000 0.952000 0.561000 1.280000 ;
        RECT 0.102000 0.952000 0.192000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 1.400000 0.080000 ;
        RECT 1.055000 -0.080000 1.161000 0.122000 ;
        RECT 1.055000 -0.080000 1.145000 0.247000 ;
        RECT 0.064000 -0.080000 0.154000 0.247000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.651000 0.689000 0.741000 0.770000 ;
        RECT 0.567000 0.164000 0.658000 0.245000 ;
        RECT 0.282000 0.689000 0.373000 0.770000 ;
        RECT 0.643000 0.689000 0.741000 0.767000 ;
        RECT 0.233000 0.689000 0.407000 0.767000 ;
        RECT 0.233000 0.700000 0.741000 0.767000 ;
        RECT 0.233000 0.177000 0.294000 0.767000 ;
        RECT 0.233000 0.177000 0.658000 0.232000 ;
        RECT 0.282000 0.177000 0.294000 0.770000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 1.262000 0.279000 1.352000 0.379000 ;
        RECT 1.262000 0.702000 1.352000 0.783000 ;
        RECT 0.567000 0.410000 0.658000 0.490000 ;
        RECT 1.140000 0.324000 1.201000 0.757000 ;
        RECT 0.597000 0.324000 0.658000 0.490000 ;
        RECT 1.140000 0.702000 1.352000 0.757000 ;
        RECT 0.597000 0.324000 1.352000 0.379000 ;
    END
END NAND3BX2

MACRO NAND3X4
    CLASS CORE ;
    FOREIGN NAND3X4 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.800000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.486000 0.426000 1.579000 0.590000 ;
        RECT 0.584000 0.411000 0.676000 0.492000 ;
        RECT 1.484000 0.426000 1.579000 0.499000 ;
        RECT 1.484000 0.302000 1.546000 0.499000 ;
        RECT 0.614000 0.302000 0.676000 0.492000 ;
        RECT 1.486000 0.302000 1.546000 0.590000 ;
        RECT 0.614000 0.302000 1.546000 0.357000 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.302000 0.494000 1.395000 0.590000 ;
        RECT 0.385000 0.514000 0.477000 0.601000 ;
        RECT 0.835000 0.417000 0.927000 0.498000 ;
        RECT 0.758000 0.418000 0.927000 0.498000 ;
        RECT 1.302000 0.418000 1.365000 0.590000 ;
        RECT 0.758000 0.418000 0.821000 0.601000 ;
        RECT 0.758000 0.418000 1.365000 0.473000 ;
        RECT 0.385000 0.546000 0.821000 0.601000 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.059000 0.439000 0.155000 0.573000 ;
        RECT 1.020000 0.527000 1.113000 0.608000 ;
        RECT 1.035000 0.527000 1.098000 0.880000 ;
        RECT 0.093000 0.439000 0.155000 0.880000 ;
        RECT 0.093000 0.825000 1.098000 0.880000 ;
        END
    END C
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 1.800000 1.280000 ;
        RECT 1.602000 0.952000 1.695000 1.280000 ;
        RECT 1.231000 0.952000 1.324000 1.280000 ;
        RECT 0.863000 0.952000 0.956000 1.280000 ;
        RECT 0.484000 0.952000 0.577000 1.280000 ;
        RECT 0.105000 0.952000 0.198000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 1.800000 0.080000 ;
        RECT 1.102000 -0.080000 1.195000 0.122000 ;
        RECT 0.063000 -0.080000 0.155000 0.247000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.218000 0.167000 0.322000 0.500000 ;
        RECT 1.620000 0.158000 1.713000 0.351000 ;
        RECT 0.224000 0.167000 0.316000 0.770000 ;
        RECT 1.560000 0.158000 1.713000 0.248000 ;
        RECT 1.417000 0.689000 1.510000 0.770000 ;
        RECT 0.224000 0.689000 0.770000 0.770000 ;
        RECT 0.218000 0.167000 0.676000 0.248000 ;
        RECT 1.645000 0.158000 1.707000 0.744000 ;
        RECT 1.417000 0.689000 1.707000 0.744000 ;
        RECT 0.218000 0.193000 1.713000 0.248000 ;
        END
    END Y
END NAND3X4

MACRO NAND3X2
    CLASS CORE ;
    FOREIGN NAND3X2 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.300000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.602000 0.300000 0.698000 0.490000 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.782000 0.433000 0.907000 0.588000 ;
        RECT 0.782000 0.493000 0.923000 0.588000 ;
        RECT 0.377000 0.514000 0.473000 0.604000 ;
        RECT 0.782000 0.433000 0.868000 0.604000 ;
        RECT 0.377000 0.549000 0.868000 0.604000 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.087000 0.460000 0.183000 0.573000 ;
        RECT 1.016000 0.573000 1.111000 0.706000 ;
        RECT 0.087000 0.439000 0.167000 0.573000 ;
        RECT 1.031000 0.573000 1.096000 0.881000 ;
        RECT 0.118000 0.460000 0.183000 0.881000 ;
        RECT 0.118000 0.826000 1.096000 0.881000 ;
        RECT 0.060000 0.439000 0.167000 0.494000 ;
        RECT 0.118000 0.439000 0.167000 0.881000 ;
        END
    END C
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 1.300000 1.280000 ;
        RECT 0.499000 0.952000 0.595000 1.280000 ;
        RECT 0.108000 0.952000 0.204000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 1.300000 0.080000 ;
        RECT 1.137000 -0.080000 1.232000 0.122000 ;
        RECT 0.068000 -0.080000 0.163000 0.122000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.691000 0.689000 0.786000 0.770000 ;
        RECT 0.602000 0.164000 0.698000 0.245000 ;
        RECT 0.300000 0.689000 0.432000 0.770000 ;
        RECT 0.682000 0.689000 0.786000 0.761000 ;
        RECT 0.248000 0.689000 0.432000 0.761000 ;
        RECT 0.300000 0.700000 0.518000 0.770000 ;
        RECT 0.248000 0.190000 0.312000 0.761000 ;
        RECT 0.248000 0.700000 0.518000 0.761000 ;
        RECT 0.248000 0.706000 0.786000 0.761000 ;
        RECT 0.248000 0.190000 0.698000 0.245000 ;
        RECT 0.300000 0.190000 0.312000 0.770000 ;
        END
    END Y
END NAND3X2

MACRO NAND3X1
    CLASS CORE ;
    FOREIGN NAND3X1 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 0.700000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.439000 0.501000 0.529000 0.582000 ;
        RECT 0.439000 0.306000 0.500000 0.582000 ;
        RECT 0.407000 0.306000 0.500000 0.361000 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.232000 0.544000 0.349000 0.676000 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.050000 0.425000 0.141000 0.590000 ;
        END
    END C
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.048000 1.078000 0.483000 1.280000 ;
        RECT 0.000000 1.120000 0.700000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 0.700000 0.080000 ;
        RECT 0.064000 -0.080000 0.154000 0.122000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.562000 0.167000 0.652000 0.307000 ;
        RECT 0.562000 0.731000 0.655000 0.812000 ;
        RECT 0.203000 0.731000 0.293000 0.812000 ;
        RECT 0.581000 0.695000 0.655000 0.812000 ;
        RECT 0.591000 0.167000 0.652000 0.812000 ;
        RECT 0.203000 0.744000 0.655000 0.799000 ;
        END
    END Y
END NAND3X1

MACRO NAND2BXL
    CLASS CORE ;
    FOREIGN NAND2BXL 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 0.700000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN AN
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.056000 0.901000 0.196000 1.033000 ;
        END
    END AN
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.232000 0.439000 0.377000 0.544000 ;
        RECT 0.212000 0.460000 0.391000 0.544000 ;
        END
    END B
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.377000 1.078000 0.636000 1.280000 ;
        RECT 0.000000 1.120000 0.700000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 0.700000 0.080000 ;
        RECT 0.207000 -0.080000 0.297000 0.122000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.557000 0.245000 0.647000 0.361000 ;
        RECT 0.398000 0.777000 0.488000 0.858000 ;
        RECT 0.601000 0.306000 0.662000 0.845000 ;
        RECT 0.407000 0.306000 0.662000 0.361000 ;
        RECT 0.398000 0.790000 0.662000 0.845000 ;
        RECT 0.601000 0.245000 0.647000 0.845000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.048000 0.740000 0.138000 0.821000 ;
        RECT 0.048000 0.274000 0.138000 0.355000 ;
        RECT 0.062000 0.668000 0.138000 0.821000 ;
        RECT 0.476000 0.613000 0.537000 0.723000 ;
        RECT 0.062000 0.274000 0.123000 0.821000 ;
        RECT 0.062000 0.668000 0.537000 0.723000 ;
    END
END NAND2BXL

MACRO NAND2BX2
    CLASS CORE ;
    FOREIGN NAND2BX2 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.100000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN AN
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.047000 0.452000 0.142000 0.627000 ;
        END
    END AN
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.853000 0.549000 0.939000 0.636000 ;
        RECT 0.372000 0.560000 0.467000 0.640000 ;
        RECT 0.372000 0.573000 0.939000 0.627000 ;
        END
    END B
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.353000 1.078000 1.050000 1.280000 ;
        RECT 0.000000 1.120000 1.100000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 1.100000 0.080000 ;
        RECT 0.233000 -0.080000 0.328000 0.122000 ;
        RECT 0.956000 -0.080000 1.050000 0.278000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.800000 0.690000 0.894000 0.771000 ;
        RECT 0.600000 0.290000 0.694000 0.371000 ;
        RECT 0.444000 0.702000 0.539000 0.783000 ;
        RECT 0.772000 0.700000 1.067000 0.770000 ;
        RECT 0.444000 0.702000 0.610000 0.770000 ;
        RECT 0.812000 0.361000 0.878000 0.457000 ;
        RECT 1.003000 0.402000 1.067000 0.770000 ;
        RECT 0.812000 0.317000 0.876000 0.457000 ;
        RECT 0.812000 0.402000 1.067000 0.457000 ;
        RECT 0.444000 0.715000 1.067000 0.770000 ;
        RECT 0.600000 0.317000 0.876000 0.371000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.050000 0.279000 0.144000 0.368000 ;
        RECT 0.639000 0.433000 0.733000 0.514000 ;
        RECT 0.050000 0.702000 0.144000 0.783000 ;
        RECT 0.049000 0.292000 0.144000 0.368000 ;
        RECT 0.208000 0.311000 0.272000 0.757000 ;
        RECT 0.049000 0.311000 0.272000 0.368000 ;
        RECT 0.272000 0.446000 0.639000 0.501000 ;
        RECT 0.050000 0.702000 0.272000 0.757000 ;
    END
END NAND2BX2

MACRO NAND2BX1
    CLASS CORE ;
    FOREIGN NAND2BX1 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 0.700000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN AN
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.056000 0.901000 0.196000 1.033000 ;
        END
    END AN
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.232000 0.439000 0.377000 0.545000 ;
        RECT 0.212000 0.461000 0.391000 0.545000 ;
        END
    END B
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.377000 1.078000 0.636000 1.280000 ;
        RECT 0.000000 1.120000 0.700000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 0.700000 0.080000 ;
        RECT 0.207000 -0.080000 0.297000 0.122000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.557000 0.289000 0.647000 0.370000 ;
        RECT 0.467000 0.300000 0.647000 0.367000 ;
        RECT 0.586000 0.289000 0.647000 0.808000 ;
        RECT 0.407000 0.306000 0.647000 0.361000 ;
        RECT 0.398000 0.754000 0.647000 0.808000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.048000 0.740000 0.138000 0.821000 ;
        RECT 0.048000 0.274000 0.138000 0.355000 ;
        RECT 0.463000 0.605000 0.524000 0.694000 ;
        RECT 0.062000 0.274000 0.123000 0.821000 ;
        RECT 0.138000 0.605000 0.524000 0.660000 ;
        RECT 0.123000 0.605000 0.463000 0.660000 ;
        RECT 0.062000 0.605000 0.138000 0.660000 ;
    END
END NAND2BX1

MACRO NAND2X4
    CLASS CORE ;
    FOREIGN NAND2X4 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.300000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.968000 0.467000 1.089000 0.573000 ;
        RECT 0.605000 0.439000 0.695000 0.521000 ;
        RECT 0.431000 0.471000 0.526000 0.552000 ;
        RECT 0.446000 0.467000 0.526000 0.552000 ;
        RECT 1.024000 0.467000 1.089000 0.652000 ;
        RECT 0.446000 0.467000 1.089000 0.521000 ;
        RECT 0.431000 0.471000 1.089000 0.521000 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.184000 0.573000 0.311000 0.662000 ;
        RECT 0.764000 0.576000 0.860000 0.657000 ;
        RECT 0.169000 0.573000 0.311000 0.654000 ;
        RECT 0.764000 0.576000 0.844000 0.662000 ;
        RECT 0.184000 0.607000 0.844000 0.662000 ;
        RECT 0.184000 0.607000 0.860000 0.657000 ;
        END
    END B
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 1.300000 1.280000 ;
        RECT 1.131000 0.871000 1.227000 1.280000 ;
        RECT 0.771000 0.871000 0.867000 1.280000 ;
        RECT 0.411000 0.871000 0.506000 1.280000 ;
        RECT 0.051000 0.871000 0.146000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 1.300000 0.080000 ;
        RECT 0.794000 -0.080000 0.889000 0.237000 ;
        RECT 0.079000 -0.080000 0.174000 0.122000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.154000 0.245000 1.261000 0.633000 ;
        RECT 0.433000 0.283000 0.529000 0.379000 ;
        RECT 1.154000 0.245000 1.249000 0.798000 ;
        RECT 0.231000 0.717000 1.249000 0.798000 ;
        RECT 0.433000 0.307000 1.261000 0.379000 ;
        END
    END Y
END NAND2X4

MACRO NAND2X2
    CLASS CORE ;
    FOREIGN NAND2X2 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 0.900000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.398000 0.400000 0.551000 0.520000 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.668000 0.558000 0.731000 0.645000 ;
        RECT 0.200000 0.573000 0.301000 0.632000 ;
        RECT 0.200000 0.577000 0.731000 0.632000 ;
        RECT 0.185000 0.573000 0.301000 0.627000 ;
        RECT 0.185000 0.577000 0.731000 0.627000 ;
        END
    END B
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.210000 1.078000 0.851000 1.280000 ;
        RECT 0.000000 1.120000 0.900000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 0.900000 0.080000 ;
        RECT 0.758000 -0.080000 0.851000 0.289000 ;
        RECT 0.049000 -0.080000 0.142000 0.122000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.409000 0.223000 0.502000 0.304000 ;
        RECT 0.779000 0.704000 0.858000 0.770000 ;
        RECT 0.795000 0.402000 0.858000 0.770000 ;
        RECT 0.618000 0.249000 0.680000 0.457000 ;
        RECT 0.599000 0.249000 0.680000 0.306000 ;
        RECT 0.618000 0.402000 0.858000 0.457000 ;
        RECT 0.409000 0.249000 0.680000 0.304000 ;
        RECT 0.251000 0.704000 0.858000 0.758000 ;
        END
    END Y
END NAND2X2

MACRO NAND2X1
    CLASS CORE ;
    FOREIGN NAND2X1 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 0.600000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.242000 0.530000 0.421000 0.633000 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.042000 0.438000 0.158000 0.598000 ;
        END
    END B
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.055000 1.078000 0.359000 1.280000 ;
        RECT 0.000000 1.120000 0.600000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 0.600000 0.080000 ;
        RECT 0.055000 -0.080000 0.158000 0.328000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.442000 0.282000 0.545000 0.367000 ;
        RECT 0.248000 0.688000 0.352000 0.769000 ;
        RECT 0.494000 0.300000 0.564000 0.743000 ;
        RECT 0.442000 0.300000 0.564000 0.367000 ;
        RECT 0.248000 0.688000 0.564000 0.743000 ;
        RECT 0.494000 0.282000 0.545000 0.743000 ;
        END
    END Y
END NAND2X1

MACRO MXI2XL
    CLASS CORE ;
    FOREIGN MXI2XL 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.300000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.128000 0.433000 1.261000 0.543000 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.411000 0.433000 0.529000 0.555000 ;
        END
    END B
    PIN S0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.198000 0.524000 0.332000 0.633000 ;
        END
    END S0
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 1.300000 1.280000 ;
        RECT 1.152000 1.064000 1.251000 1.280000 ;
        RECT 0.304000 0.941000 0.400000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 1.300000 0.080000 ;
        RECT 1.151000 -0.080000 1.247000 0.122000 ;
        RECT 0.308000 -0.080000 0.404000 0.347000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.764000 0.573000 0.868000 0.819000 ;
        RECT 0.748000 0.738000 0.868000 0.819000 ;
        RECT 0.748000 0.281000 0.844000 0.362000 ;
        RECT 0.764000 0.281000 0.829000 0.819000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.049000 0.779000 0.152000 0.870000 ;
        RECT 0.974000 0.738000 1.069000 0.819000 ;
        RECT 0.962000 0.279000 1.058000 0.360000 ;
        RECT 0.590000 0.930000 0.698000 1.011000 ;
        RECT 0.535000 0.281000 0.677000 0.362000 ;
        RECT 0.529000 0.679000 0.677000 0.760000 ;
        RECT 0.049000 0.281000 0.163000 0.362000 ;
        RECT 0.975000 0.279000 1.040000 0.819000 ;
        RECT 0.612000 0.281000 0.677000 0.760000 ;
        RECT 0.049000 0.281000 0.114000 0.870000 ;
        RECT 0.590000 0.815000 0.654000 1.011000 ;
        RECT 0.049000 0.815000 0.654000 0.870000 ;
    END
END MXI2XL

MACRO MX2XL
    CLASS CORE ;
    FOREIGN MX2XL 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.400000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.000000 0.419000 1.188000 0.513000 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.387000 0.654000 0.488000 0.767000 ;
        RECT 0.292000 0.619000 0.387000 0.730000 ;
        RECT 0.292000 0.654000 0.488000 0.730000 ;
        END
    END B
    PIN S0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.037000 0.958000 0.188000 1.048000 ;
        END
    END S0
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 1.400000 1.280000 ;
        RECT 1.050000 1.078000 1.140000 1.280000 ;
        RECT 0.251000 0.838000 0.341000 1.280000 ;
        RECT 0.239000 0.800000 0.326000 0.889000 ;
        RECT 0.251000 0.800000 0.326000 1.280000 ;
        RECT 0.239000 0.838000 0.341000 0.889000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 1.400000 0.080000 ;
        RECT 1.049000 -0.080000 1.139000 0.122000 ;
        RECT 0.264000 -0.080000 0.349000 0.342000 ;
        RECT 0.261000 0.291000 0.351000 0.342000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.248000 0.268000 1.363000 0.361000 ;
        RECT 1.282000 0.761000 1.363000 0.845000 ;
        RECT 1.198000 0.764000 1.363000 0.845000 ;
        RECT 1.302000 0.268000 1.363000 0.845000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.671000 0.789000 0.793000 0.882000 ;
        RECT 0.460000 0.507000 0.546000 0.599000 ;
        RECT 0.862000 0.276000 0.944000 0.358000 ;
        RECT 1.103000 0.579000 1.193000 0.660000 ;
        RECT 0.473000 0.275000 0.563000 0.356000 ;
        RECT 0.048000 0.788000 0.138000 0.869000 ;
        RECT 0.048000 0.276000 0.138000 0.357000 ;
        RECT 1.103000 0.579000 1.179000 0.676000 ;
        RECT 1.035000 0.621000 1.096000 0.968000 ;
        RECT 0.862000 0.276000 0.923000 0.819000 ;
        RECT 0.732000 0.280000 0.793000 0.968000 ;
        RECT 0.610000 0.393000 0.671000 0.720000 ;
        RECT 0.549000 0.665000 0.610000 0.906000 ;
        RECT 0.502000 0.275000 0.563000 0.448000 ;
        RECT 0.062000 0.276000 0.123000 0.869000 ;
        RECT 1.035000 0.621000 1.179000 0.676000 ;
        RECT 0.732000 0.913000 1.096000 0.968000 ;
        RECT 0.664000 0.280000 0.793000 0.335000 ;
        RECT 0.549000 0.665000 0.671000 0.720000 ;
        RECT 0.502000 0.393000 0.671000 0.448000 ;
        RECT 0.440000 0.851000 0.610000 0.906000 ;
        RECT 0.138000 0.507000 0.546000 0.562000 ;
        RECT 0.123000 0.507000 0.460000 0.562000 ;
        RECT 0.062000 0.507000 0.440000 0.562000 ;
    END
END MX2XL

MACRO INVXL
    CLASS CORE ;
    FOREIGN INVXL 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 0.400000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.042000 0.433000 0.158000 0.598000 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 0.400000 1.280000 ;
        RECT 0.155000 0.925000 0.258000 1.280000 ;
        RECT 0.083000 0.925000 0.329000 0.975000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.055000 -0.080000 0.300000 0.122000 ;
        RECT 0.000000 -0.080000 0.400000 0.080000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.242000 0.567000 0.358000 0.768000 ;
        RECT 0.236000 0.321000 0.339000 0.439000 ;
        RECT 0.242000 0.321000 0.312000 0.768000 ;
        END
    END Y
END INVXL

MACRO INVX8
    CLASS CORE ;
    FOREIGN INVX8 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.100000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.150000 0.487000 0.376000 0.633000 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.828000 1.078000 1.050000 1.280000 ;
        RECT 0.000000 1.120000 1.100000 1.280000 ;
        RECT 0.828000 0.917000 0.922000 1.280000 ;
        RECT 0.438000 0.917000 0.532000 1.280000 ;
        RECT 0.050000 0.917000 0.144000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.818000 -0.080000 1.043000 0.122000 ;
        RECT 0.000000 -0.080000 1.100000 0.080000 ;
        RECT 0.061000 -0.080000 0.156000 0.122000 ;
        RECT 0.439000 -0.080000 0.533000 0.214000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.610000 0.419000 1.040000 0.767000 ;
        RECT 0.610000 0.361000 0.878000 0.767000 ;
        RECT 0.610000 0.361000 0.857000 0.780000 ;
        RECT 0.610000 0.307000 0.811000 0.812000 ;
        RECT 0.589000 0.307000 0.811000 0.433000 ;
        RECT 0.217000 0.698000 0.811000 0.812000 ;
        RECT 0.217000 0.307000 0.811000 0.421000 ;
        RECT 0.217000 0.698000 0.857000 0.780000 ;
        RECT 0.589000 0.361000 0.878000 0.433000 ;
        RECT 0.217000 0.698000 1.040000 0.767000 ;
        RECT 0.217000 0.361000 0.878000 0.421000 ;
        END
    END Y
END INVX8

MACRO INVX4
    CLASS CORE ;
    FOREIGN INVX4 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 0.700000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.037000 0.446000 0.138000 0.633000 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 0.700000 1.280000 ;
        RECT 0.452000 0.720000 0.542000 1.280000 ;
        RECT 0.048000 0.720000 0.138000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 0.700000 0.080000 ;
        RECT 0.452000 -0.080000 0.542000 0.372000 ;
        RECT 0.048000 -0.080000 0.138000 0.372000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.212000 0.433000 0.341000 0.767000 ;
        RECT 0.251000 0.194000 0.341000 1.010000 ;
        END
    END Y
END INVX4

MACRO INVX3
    CLASS CORE ;
    FOREIGN INVX3 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 0.700000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.037000 0.493000 0.266000 0.633000 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 0.700000 1.280000 ;
        RECT 0.251000 1.078000 0.341000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 0.700000 0.080000 ;
        RECT 0.251000 -0.080000 0.341000 0.122000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.387000 0.700000 0.489000 0.900000 ;
        RECT 0.399000 0.295000 0.489000 0.913000 ;
        RECT 0.049000 0.720000 0.139000 0.913000 ;
        RECT 0.049000 0.215000 0.139000 0.408000 ;
        RECT 0.049000 0.773000 0.489000 0.854000 ;
        RECT 0.049000 0.295000 0.489000 0.376000 ;
        END
    END Y
END INVX3

MACRO INVX2
    CLASS CORE ;
    FOREIGN INVX2 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 0.600000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.150000 0.433000 0.395000 0.574000 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 0.600000 1.280000 ;
        RECT 0.394000 1.078000 0.497000 1.280000 ;
        RECT 0.395000 1.064000 0.495000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 0.600000 0.080000 ;
        RECT 0.164000 -0.080000 0.267000 0.361000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.442000 0.183000 0.558000 0.376000 ;
        RECT 0.224000 0.661000 0.327000 0.854000 ;
        RECT 0.465000 0.627000 0.558000 0.715000 ;
        RECT 0.488000 0.183000 0.558000 0.715000 ;
        RECT 0.224000 0.661000 0.558000 0.715000 ;
        END
    END Y
END INVX2

MACRO INVX1
    CLASS CORE ;
    FOREIGN INVX1 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 0.400000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.042000 0.433000 0.173000 0.568000 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 0.400000 1.280000 ;
        RECT 0.055000 1.078000 0.158000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 0.400000 0.080000 ;
        RECT 0.055000 -0.080000 0.158000 0.122000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.242000 0.564000 0.358000 0.848000 ;
        RECT 0.253000 0.321000 0.323000 0.848000 ;
        END
    END Y
END INVX1

MACRO INVX12
    CLASS CORE ;
    FOREIGN INVX12 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 2.300000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.139000 0.507000 0.231000 0.588000 ;
        RECT 0.058000 0.533000 0.119000 0.627000 ;
        RECT 0.058000 0.533000 0.231000 0.588000 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 2.300000 1.280000 ;
        RECT 1.017000 1.065000 1.110000 1.280000 ;
        RECT 2.161000 0.989000 2.252000 1.280000 ;
        RECT 1.777000 0.989000 1.868000 1.280000 ;
        RECT 1.393000 0.989000 1.484000 1.280000 ;
        RECT 0.268000 1.078000 0.359000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 2.300000 0.080000 ;
        RECT 2.158000 -0.080000 2.249000 0.199000 ;
        RECT 1.777000 -0.080000 1.868000 0.199000 ;
        RECT 1.393000 -0.080000 1.484000 0.199000 ;
        RECT 0.654000 -0.080000 0.745000 0.122000 ;
        RECT 0.283000 -0.080000 0.374000 0.237000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.827000 0.286000 2.242000 0.914000 ;
        RECT 1.807000 0.626000 2.242000 0.914000 ;
        RECT 1.154000 0.676000 2.242000 0.914000 ;
        RECT 1.155000 0.286000 2.242000 0.448000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.470000 0.686000 0.562000 0.888000 ;
        RECT 0.855000 0.521000 1.745000 0.602000 ;
        RECT 0.855000 0.338000 0.936000 0.767000 ;
        RECT 0.470000 0.686000 0.936000 0.767000 ;
        RECT 0.470000 0.338000 0.936000 0.419000 ;
        RECT 0.318000 0.500000 0.713000 0.581000 ;
        RECT 0.054000 0.343000 0.145000 0.424000 ;
        RECT 0.048000 0.689000 0.139000 0.770000 ;
        RECT 0.318000 0.343000 0.379000 0.770000 ;
        RECT 0.054000 0.343000 0.379000 0.398000 ;
        RECT 0.048000 0.715000 0.379000 0.770000 ;
    END
END INVX12

MACRO DLY4X1
    CLASS CORE ;
    FOREIGN DLY4X1 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.300000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.129000 0.860000 0.225000 0.940000 ;
        RECT 0.129000 0.860000 0.311000 0.927000 ;
        RECT 0.246000 0.839000 0.311000 0.927000 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 1.300000 1.280000 ;
        RECT 0.996000 1.078000 1.092000 1.280000 ;
        RECT 0.242000 1.078000 0.338000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 1.300000 0.080000 ;
        RECT 0.996000 -0.080000 1.092000 0.122000 ;
        RECT 0.310000 -0.080000 0.405000 0.122000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.154000 0.738000 1.249000 0.819000 ;
        RECT 1.154000 0.312000 1.249000 0.393000 ;
        RECT 1.175000 0.706000 1.249000 0.819000 ;
        RECT 1.185000 0.312000 1.249000 0.819000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.926000 0.486000 1.119000 0.567000 ;
        RECT 0.650000 0.486000 0.861000 0.567000 ;
        RECT 0.619000 0.652000 0.715000 0.733000 ;
        RECT 0.619000 0.336000 0.715000 0.417000 ;
        RECT 0.619000 0.170000 0.715000 0.251000 ;
        RECT 0.588000 0.840000 0.684000 0.921000 ;
        RECT 0.082000 0.517000 0.484000 0.598000 ;
        RECT 0.051000 0.652000 0.146000 0.733000 ;
        RECT 0.051000 0.336000 0.146000 0.417000 ;
        RECT 0.650000 0.336000 0.715000 0.733000 ;
        RECT 0.926000 0.196000 0.990000 0.895000 ;
        RECT 0.082000 0.336000 0.146000 0.733000 ;
        RECT 0.619000 0.196000 0.990000 0.251000 ;
        RECT 0.588000 0.840000 0.990000 0.895000 ;
    END
END DLY4X1

MACRO DLY3X1
    CLASS CORE ;
    FOREIGN DLY3X1 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.300000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.129000 0.860000 0.225000 0.940000 ;
        RECT 0.129000 0.860000 0.311000 0.927000 ;
        RECT 0.246000 0.839000 0.311000 0.927000 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 1.300000 1.280000 ;
        RECT 0.937000 1.078000 1.035000 1.280000 ;
        RECT 0.259000 1.078000 0.355000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 1.300000 0.080000 ;
        RECT 0.937000 -0.080000 1.033000 0.122000 ;
        RECT 0.259000 -0.080000 0.355000 0.122000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.154000 0.738000 1.249000 0.819000 ;
        RECT 1.154000 0.312000 1.249000 0.393000 ;
        RECT 1.175000 0.706000 1.249000 0.819000 ;
        RECT 1.185000 0.312000 1.249000 0.819000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.895000 0.486000 1.113000 0.567000 ;
        RECT 0.616000 0.486000 0.830000 0.567000 ;
        RECT 0.588000 0.840000 0.684000 0.921000 ;
        RECT 0.588000 0.170000 0.684000 0.251000 ;
        RECT 0.585000 0.652000 0.681000 0.733000 ;
        RECT 0.585000 0.336000 0.681000 0.417000 ;
        RECT 0.082000 0.517000 0.501000 0.598000 ;
        RECT 0.051000 0.652000 0.146000 0.733000 ;
        RECT 0.051000 0.336000 0.146000 0.417000 ;
        RECT 0.895000 0.196000 0.960000 0.895000 ;
        RECT 0.616000 0.336000 0.681000 0.733000 ;
        RECT 0.082000 0.336000 0.146000 0.733000 ;
        RECT 0.588000 0.840000 0.960000 0.895000 ;
        RECT 0.588000 0.196000 0.960000 0.251000 ;
    END
END DLY3X1

MACRO DLY2X1
    CLASS CORE ;
    FOREIGN DLY2X1 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.100000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.128000 0.860000 0.222000 0.940000 ;
        RECT 0.128000 0.860000 0.307000 0.927000 ;
        RECT 0.243000 0.839000 0.307000 0.927000 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 1.100000 1.280000 ;
        RECT 0.800000 1.078000 0.894000 1.280000 ;
        RECT 0.256000 1.078000 0.350000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 1.100000 0.080000 ;
        RECT 0.800000 -0.080000 0.894000 0.122000 ;
        RECT 0.256000 -0.080000 0.350000 0.122000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.956000 0.738000 1.050000 0.819000 ;
        RECT 0.956000 0.312000 1.050000 0.393000 ;
        RECT 0.976000 0.706000 1.050000 0.819000 ;
        RECT 0.986000 0.312000 1.050000 0.819000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.828000 0.486000 0.921000 0.567000 ;
        RECT 0.558000 0.486000 0.750000 0.567000 ;
        RECT 0.528000 0.840000 0.622000 0.921000 ;
        RECT 0.528000 0.652000 0.622000 0.733000 ;
        RECT 0.528000 0.336000 0.622000 0.417000 ;
        RECT 0.528000 0.170000 0.622000 0.251000 ;
        RECT 0.081000 0.517000 0.478000 0.598000 ;
        RECT 0.050000 0.652000 0.144000 0.733000 ;
        RECT 0.050000 0.336000 0.144000 0.417000 ;
        RECT 0.828000 0.196000 0.892000 0.895000 ;
        RECT 0.558000 0.336000 0.622000 0.733000 ;
        RECT 0.081000 0.336000 0.144000 0.733000 ;
        RECT 0.528000 0.840000 0.892000 0.895000 ;
        RECT 0.528000 0.196000 0.892000 0.251000 ;
    END
END DLY2X1

MACRO DLY1X1
    CLASS CORE ;
    FOREIGN DLY1X1 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.100000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.125000 0.826000 0.219000 0.907000 ;
        RECT 0.125000 0.826000 0.243000 0.900000 ;
        RECT 0.125000 0.833000 0.328000 0.900000 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 1.100000 1.280000 ;
        RECT 0.744000 1.078000 0.839000 1.280000 ;
        RECT 0.300000 1.078000 0.394000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 1.100000 0.080000 ;
        RECT 0.744000 -0.080000 0.839000 0.122000 ;
        RECT 0.300000 -0.080000 0.394000 0.122000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.956000 0.760000 1.050000 0.857000 ;
        RECT 0.956000 0.243000 1.050000 0.324000 ;
        RECT 0.976000 0.243000 1.040000 0.857000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.758000 0.486000 0.892000 0.567000 ;
        RECT 0.553000 0.486000 0.694000 0.567000 ;
        RECT 0.522000 0.840000 0.617000 0.921000 ;
        RECT 0.522000 0.652000 0.617000 0.733000 ;
        RECT 0.522000 0.336000 0.617000 0.417000 ;
        RECT 0.081000 0.517000 0.472000 0.598000 ;
        RECT 0.050000 0.652000 0.144000 0.733000 ;
        RECT 0.050000 0.336000 0.144000 0.417000 ;
        RECT 0.522000 0.170000 0.617000 0.246000 ;
        RECT 0.758000 0.192000 0.822000 0.895000 ;
        RECT 0.553000 0.336000 0.617000 0.733000 ;
        RECT 0.081000 0.336000 0.144000 0.733000 ;
        RECT 0.522000 0.840000 0.822000 0.895000 ;
        RECT 0.522000 0.192000 0.822000 0.246000 ;
    END
END DLY1X1

MACRO BUFX8
    CLASS CORE ;
    FOREIGN BUFX8 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.600000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.154000 0.474000 0.372000 0.555000 ;
        RECT 0.236000 0.439000 0.298000 0.555000 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 1.600000 1.280000 ;
        RECT 1.104000 0.877000 1.196000 1.280000 ;
        RECT 0.070000 0.897000 0.162000 1.280000 ;
        RECT 0.760000 0.877000 0.851000 1.280000 ;
        RECT 0.415000 0.897000 0.506000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 1.600000 0.080000 ;
        RECT 1.126000 -0.080000 1.218000 0.211000 ;
        RECT 0.781000 -0.080000 0.873000 0.211000 ;
        RECT 0.436000 -0.080000 0.528000 0.198000 ;
        RECT 0.048000 -0.080000 0.140000 0.211000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.947000 0.433000 1.364000 0.767000 ;
        RECT 0.947000 0.433000 1.220000 0.774000 ;
        RECT 0.947000 0.307000 1.131000 0.774000 ;
        RECT 0.927000 0.626000 1.220000 0.774000 ;
        RECT 0.927000 0.626000 1.364000 0.767000 ;
        RECT 0.927000 0.307000 1.131000 0.440000 ;
        RECT 0.609000 0.307000 1.131000 0.421000 ;
        RECT 0.587000 0.660000 1.220000 0.774000 ;
        RECT 0.587000 0.660000 1.364000 0.767000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.434000 0.274000 0.525000 0.738000 ;
        RECT 0.434000 0.519000 0.865000 0.600000 ;
        RECT 0.242000 0.657000 0.525000 0.738000 ;
        RECT 0.242000 0.274000 0.525000 0.355000 ;
    END
END BUFX8

MACRO BUFX4
    CLASS CORE ;
    FOREIGN BUFX4 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 0.900000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.038000 0.433000 0.218000 0.570000 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 0.900000 1.280000 ;
        RECT 0.671000 0.953000 0.764000 1.280000 ;
        RECT 0.256000 0.953000 0.349000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 0.900000 0.080000 ;
        RECT 0.671000 -0.080000 0.764000 0.122000 ;
        RECT 0.256000 -0.080000 0.349000 0.122000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.464000 0.652000 0.600000 0.767000 ;
        RECT 0.464000 0.300000 0.682000 0.412000 ;
        RECT 0.578000 0.300000 0.682000 0.733000 ;
        RECT 0.464000 0.652000 0.556000 0.957000 ;
        RECT 0.464000 0.219000 0.556000 0.412000 ;
        RECT 0.464000 0.652000 0.682000 0.733000 ;
        RECT 0.578000 0.300000 0.600000 0.767000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.284000 0.477000 0.515000 0.585000 ;
        RECT 0.049000 0.652000 0.142000 0.957000 ;
        RECT 0.049000 0.186000 0.142000 0.379000 ;
        RECT 0.284000 0.298000 0.376000 0.733000 ;
        RECT 0.049000 0.652000 0.376000 0.733000 ;
        RECT 0.049000 0.298000 0.376000 0.379000 ;
    END
END BUFX4

MACRO BUFX3
    CLASS CORE ;
    FOREIGN BUFX3 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 0.700000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.037000 0.433000 0.147000 0.562000 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 0.700000 1.280000 ;
        RECT 0.196000 1.078000 0.286000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 0.700000 0.080000 ;
        RECT 0.557000 -0.080000 0.647000 0.122000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.387000 0.433000 0.488000 0.633000 ;
        RECT 0.398000 0.433000 0.488000 0.752000 ;
        RECT 0.408000 0.287000 0.498000 0.368000 ;
        RECT 0.408000 0.287000 0.469000 0.752000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.235000 0.470000 0.325000 0.551000 ;
        RECT 0.048000 0.696000 0.138000 0.777000 ;
        RECT 0.048000 0.244000 0.138000 0.325000 ;
        RECT 0.235000 0.270000 0.296000 0.751000 ;
        RECT 0.048000 0.696000 0.296000 0.751000 ;
        RECT 0.048000 0.270000 0.296000 0.325000 ;
    END
END BUFX3

MACRO BUFX2
    CLASS CORE ;
    FOREIGN BUFX2 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 0.700000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.037000 0.418000 0.236000 0.538000 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 0.700000 1.280000 ;
        RECT 0.223000 1.078000 0.313000 1.280000 ;
        RECT 0.237000 1.065000 0.298000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 0.700000 0.080000 ;
        RECT 0.233000 -0.080000 0.323000 0.122000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.435000 0.331000 0.525000 0.412000 ;
        RECT 0.424000 0.655000 0.514000 0.736000 ;
        RECT 0.562000 0.357000 0.623000 0.710000 ;
        RECT 0.562000 0.439000 0.643000 0.494000 ;
        RECT 0.435000 0.357000 0.623000 0.412000 ;
        RECT 0.424000 0.655000 0.623000 0.710000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.302000 0.490000 0.430000 0.571000 ;
        RECT 0.074000 0.657000 0.164000 0.738000 ;
        RECT 0.074000 0.275000 0.164000 0.356000 ;
        RECT 0.302000 0.301000 0.363000 0.712000 ;
        RECT 0.074000 0.657000 0.363000 0.712000 ;
        RECT 0.074000 0.301000 0.363000 0.356000 ;
    END
END BUFX2

MACRO BUFX20
    CLASS CORE ;
    FOREIGN BUFX20 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 2.800000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.199000 0.474000 0.663000 0.555000 ;
        RECT 0.407000 0.439000 0.468000 0.555000 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 2.800000 1.280000 ;
        RECT 2.434000 1.078000 2.524000 1.280000 ;
        RECT 2.084000 0.989000 2.174000 1.280000 ;
        RECT 1.745000 0.989000 1.835000 1.280000 ;
        RECT 1.405000 0.972000 1.495000 1.280000 ;
        RECT 1.066000 0.972000 1.156000 1.280000 ;
        RECT 0.727000 0.873000 0.817000 1.280000 ;
        RECT 0.387000 0.873000 0.477000 1.280000 ;
        RECT 0.048000 0.873000 0.138000 1.280000 ;
        RECT 2.449000 1.065000 2.510000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 2.800000 0.080000 ;
        RECT 2.445000 -0.080000 2.535000 0.122000 ;
        RECT 2.095000 -0.080000 2.185000 0.198000 ;
        RECT 1.755000 -0.080000 1.845000 0.198000 ;
        RECT 1.416000 -0.080000 1.506000 0.198000 ;
        RECT 1.077000 -0.080000 1.167000 0.198000 ;
        RECT 0.737000 -0.080000 0.827000 0.215000 ;
        RECT 0.387000 -0.080000 0.477000 0.234000 ;
        RECT 0.048000 -0.080000 0.138000 0.234000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 2.332000 0.268000 2.743000 0.914000 ;
        RECT 2.312000 0.683000 2.743000 0.839000 ;
        RECT 0.907000 0.268000 2.743000 0.408000 ;
        RECT 0.896000 0.699000 2.743000 0.839000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.744000 0.320000 0.834000 0.757000 ;
        RECT 0.744000 0.513000 2.190000 0.594000 ;
        RECT 0.557000 0.320000 0.834000 0.401000 ;
        RECT 0.217000 0.676000 0.834000 0.757000 ;
        RECT 0.217000 0.320000 0.308000 0.401000 ;
        RECT 0.217000 0.320000 0.834000 0.375000 ;
    END
END BUFX20

MACRO BUFX16
    CLASS CORE ;
    FOREIGN BUFX16 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 2.300000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.155000 0.521000 0.547000 0.602000 ;
        RECT 0.411000 0.521000 0.473000 0.627000 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 2.300000 1.280000 ;
        RECT 1.431000 0.972000 1.523000 1.280000 ;
        RECT 0.391000 0.823000 0.483000 1.280000 ;
        RECT 2.161000 1.078000 2.252000 1.280000 ;
        RECT 1.796000 1.078000 1.887000 1.280000 ;
        RECT 1.088000 0.972000 1.179000 1.280000 ;
        RECT 0.745000 0.972000 0.836000 1.280000 ;
        RECT 0.048000 0.823000 0.139000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 2.300000 0.080000 ;
        RECT 1.978000 -0.080000 2.069000 0.122000 ;
        RECT 1.614000 -0.080000 1.705000 0.198000 ;
        RECT 1.260000 -0.080000 1.351000 0.198000 ;
        RECT 0.917000 -0.080000 1.008000 0.198000 ;
        RECT 0.563000 -0.080000 0.654000 0.216000 ;
        RECT 0.220000 -0.080000 0.311000 0.215000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.827000 0.268000 2.242000 0.914000 ;
        RECT 1.807000 0.675000 2.242000 0.839000 ;
        RECT 0.917000 0.699000 2.242000 0.839000 ;
        RECT 0.745000 0.268000 2.242000 0.408000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.563000 0.657000 0.672000 0.743000 ;
        RECT 0.220000 0.657000 0.311000 0.743000 ;
        RECT 0.610000 0.513000 1.745000 0.594000 ;
        RECT 0.048000 0.335000 0.672000 0.415000 ;
        RECT 0.610000 0.335000 0.672000 0.743000 ;
        RECT 0.220000 0.688000 0.672000 0.743000 ;
    END
END BUFX16

MACRO BUFX12
    CLASS CORE ;
    FOREIGN BUFX12 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.800000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.194000 0.474000 0.554000 0.555000 ;
        RECT 0.239000 0.439000 0.301000 0.555000 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 1.800000 1.280000 ;
        RECT 1.658000 0.972000 1.751000 1.280000 ;
        RECT 0.922000 0.972000 1.015000 1.280000 ;
        RECT 1.285000 0.972000 1.377000 1.280000 ;
        RECT 0.573000 0.897000 0.665000 1.280000 ;
        RECT 0.224000 0.897000 0.316000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 1.800000 0.080000 ;
        RECT 1.642000 -0.080000 1.735000 0.211000 ;
        RECT 1.293000 -0.080000 1.385000 0.211000 ;
        RECT 0.944000 -0.080000 1.036000 0.215000 ;
        RECT 0.595000 -0.080000 0.687000 0.215000 ;
        RECT 0.235000 -0.080000 0.327000 0.122000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.319000 0.300000 1.741000 0.767000 ;
        RECT 1.298000 0.626000 1.741000 0.757000 ;
        RECT 1.298000 0.321000 1.741000 0.440000 ;
        RECT 0.769000 0.321000 1.741000 0.402000 ;
        RECT 0.747000 0.676000 1.741000 0.757000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.622000 0.519000 1.193000 0.600000 ;
        RECT 0.420000 0.319000 0.513000 0.400000 ;
        RECT 0.398000 0.657000 0.491000 0.738000 ;
        RECT 0.049000 0.657000 0.142000 0.738000 ;
        RECT 0.622000 0.345000 0.685000 0.712000 ;
        RECT 0.079000 0.319000 0.142000 0.389000 ;
        RECT 0.420000 0.345000 0.685000 0.400000 ;
        RECT 0.079000 0.319000 0.513000 0.374000 ;
        RECT 0.049000 0.657000 0.685000 0.712000 ;
        RECT 0.049000 0.335000 0.142000 0.389000 ;
    END
END BUFX12

MACRO AOI22XL
    CLASS CORE ;
    FOREIGN AOI22XL 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 0.900000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.481000 0.412000 0.601000 0.500000 ;
        RECT 0.417000 0.425000 0.603000 0.500000 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.567000 0.562000 0.716000 0.652000 ;
        RECT 0.567000 0.571000 0.731000 0.652000 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.325000 0.560000 0.417000 0.649000 ;
        RECT 0.218000 0.567000 0.417000 0.649000 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.038000 0.396000 0.169000 0.511000 ;
        END
    END B1
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 0.900000 1.280000 ;
        RECT 0.063000 1.078000 0.176000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 0.900000 0.080000 ;
        RECT 0.747000 -0.080000 0.840000 0.122000 ;
        RECT 0.049000 -0.080000 0.142000 0.122000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.573000 0.748000 0.665000 0.829000 ;
        RECT 0.409000 0.269000 0.502000 0.350000 ;
        RECT 0.779000 0.282000 0.862000 0.361000 ;
        RECT 0.799000 0.282000 0.862000 0.815000 ;
        RECT 0.409000 0.282000 0.862000 0.337000 ;
        RECT 0.573000 0.761000 0.862000 0.815000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.049000 0.749000 0.142000 0.830000 ;
        RECT 0.390000 0.762000 0.453000 1.049000 ;
        RECT 0.390000 0.994000 0.821000 1.049000 ;
        RECT 0.142000 0.762000 0.390000 0.817000 ;
    END
END AOI22XL

MACRO AOI22X4
    CLASS CORE ;
    FOREIGN AOI22X4 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 2.500000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 2.043000 0.504000 2.105000 0.627000 ;
        RECT 1.370000 0.573000 2.105000 0.627000 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.185000 0.439000 1.247000 0.654000 ;
        RECT 1.185000 0.439000 1.288000 0.500000 ;
        RECT 1.185000 0.439000 1.872000 0.494000 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.594000 0.573000 0.656000 0.642000 ;
        RECT 0.114000 0.587000 0.770000 0.642000 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.004000 0.438000 1.066000 0.494000 ;
        RECT 1.004000 0.438000 1.081000 0.493000 ;
        RECT 0.237000 0.439000 1.066000 0.494000 ;
        RECT 0.237000 0.439000 1.081000 0.493000 ;
        END
    END B1
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 2.500000 1.280000 ;
        RECT 0.568000 0.980000 0.660000 1.280000 ;
        RECT 0.222000 0.980000 0.314000 1.280000 ;
        RECT 0.915000 0.980000 1.006000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 2.500000 0.080000 ;
        RECT 1.780000 -0.080000 1.872000 0.203000 ;
        RECT 1.088000 -0.080000 1.180000 0.203000 ;
        RECT 0.395000 -0.080000 0.487000 0.203000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 2.181000 0.439000 2.346000 0.633000 ;
        RECT 2.181000 0.300000 2.284000 0.633000 ;
        RECT 1.939000 0.930000 2.024000 1.033000 ;
        RECT 2.181000 0.287000 2.263000 0.633000 ;
        RECT 1.905000 0.967000 2.024000 1.033000 ;
        RECT 2.284000 0.439000 2.346000 0.985000 ;
        RECT 1.939000 0.930000 2.346000 0.985000 ;
        RECT 0.049000 0.287000 2.263000 0.342000 ;
        RECT 1.261000 0.979000 2.024000 1.033000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.049000 0.737000 2.219000 0.792000 ;
    END
END AOI22X4

MACRO AOI22X2
    CLASS CORE ;
    FOREIGN AOI22X2 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.600000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.061000 0.567000 1.207000 0.661000 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.356000 0.438000 1.418000 0.551000 ;
        RECT 0.882000 0.438000 0.944000 0.664000 ;
        RECT 0.882000 0.438000 1.009000 0.494000 ;
        RECT 0.882000 0.438000 1.418000 0.493000 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.329000 0.573000 0.475000 0.663000 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.185000 0.439000 0.298000 0.511000 ;
        RECT 0.113000 0.493000 0.246000 0.562000 ;
        RECT 0.653000 0.456000 0.715000 0.575000 ;
        RECT 0.185000 0.439000 0.246000 0.562000 ;
        RECT 0.185000 0.456000 0.715000 0.511000 ;
        END
    END B1
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 1.600000 1.280000 ;
        RECT 0.566000 0.888000 0.657000 1.280000 ;
        RECT 0.221000 0.888000 0.312000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 1.600000 0.080000 ;
        RECT 1.352000 -0.080000 1.444000 0.122000 ;
        RECT 0.695000 -0.080000 0.787000 0.122000 ;
        RECT 0.048000 -0.080000 0.140000 0.305000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.302000 0.706000 1.368000 0.789000 ;
        RECT 1.480000 0.321000 1.542000 0.761000 ;
        RECT 1.302000 0.706000 1.542000 0.761000 ;
        RECT 0.393000 0.321000 1.542000 0.376000 ;
        RECT 0.932000 0.735000 1.368000 0.789000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.753000 0.732000 0.815000 0.940000 ;
        RECT 0.048000 0.732000 0.830000 0.787000 ;
        RECT 0.753000 0.886000 1.541000 0.940000 ;
    END
END AOI22X2

MACRO AOI22X1
    CLASS CORE ;
    FOREIGN AOI22X1 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 0.900000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.499000 0.394000 0.592000 0.475000 ;
        RECT 0.419000 0.407000 0.592000 0.475000 ;
        RECT 0.419000 0.407000 0.481000 0.494000 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.577000 0.538000 0.731000 0.633000 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.239000 0.567000 0.415000 0.663000 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.052000 0.421000 0.145000 0.589000 ;
        END
    END B1
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 0.900000 1.280000 ;
        RECT 0.229000 1.078000 0.322000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 0.900000 0.080000 ;
        RECT 0.758000 -0.080000 0.851000 0.122000 ;
        RECT 0.049000 -0.080000 0.142000 0.330000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.779000 0.265000 0.862000 0.361000 ;
        RECT 0.584000 0.699000 0.676000 0.780000 ;
        RECT 0.398000 0.252000 0.491000 0.333000 ;
        RECT 0.799000 0.265000 0.862000 0.754000 ;
        RECT 0.584000 0.699000 0.862000 0.754000 ;
        RECT 0.398000 0.265000 0.862000 0.320000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.049000 0.726000 0.142000 0.933000 ;
        RECT 0.758000 0.854000 0.851000 0.935000 ;
        RECT 0.409000 0.865000 0.502000 0.946000 ;
        RECT 0.409000 0.880000 0.851000 0.935000 ;
        RECT 0.049000 0.879000 0.502000 0.933000 ;
        RECT 0.049000 0.880000 0.851000 0.933000 ;
    END
END AOI22X1

MACRO AOI222X4
    CLASS CORE ;
    FOREIGN AOI222X4 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 2.100000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.912000 0.398000 1.013000 0.556000 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.094000 0.524000 1.188000 0.686000 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.737000 0.505000 0.838000 0.677000 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.407000 0.573000 0.642000 0.627000 ;
        END
    END B1
    PIN C0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.231000 0.382000 0.414000 0.494000 ;
        END
    END C0
    PIN C1
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.037000 0.433000 0.138000 0.624000 ;
        END
    END C1
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 2.100000 1.280000 ;
        RECT 1.893000 0.982000 1.983000 1.280000 ;
        RECT 1.554000 0.908000 1.644000 1.280000 ;
        RECT 0.345000 1.078000 0.435000 1.280000 ;
        RECT 0.048000 1.078000 0.138000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 2.100000 0.080000 ;
        RECT 0.048000 -0.080000 0.180000 0.083000 ;
        RECT 1.893000 -0.080000 1.983000 0.212000 ;
        RECT 1.543000 -0.080000 1.633000 0.212000 ;
        RECT 1.167000 -0.080000 1.257000 0.122000 ;
        RECT 0.573000 -0.080000 0.663000 0.122000 ;
        RECT 0.048000 -0.080000 0.138000 0.275000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.787000 0.567000 1.888000 0.900000 ;
        RECT 1.787000 0.336000 1.875000 0.440000 ;
        RECT 1.723000 0.661000 1.888000 0.742000 ;
        RECT 1.814000 0.336000 1.875000 0.900000 ;
        RECT 1.723000 0.336000 1.875000 0.390000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.870000 0.236000 0.963000 0.320000 ;
        RECT 1.534000 0.287000 1.595000 0.705000 ;
        RECT 1.377000 0.650000 1.438000 0.740000 ;
        RECT 1.249000 0.404000 1.310000 0.833000 ;
        RECT 1.078000 0.265000 1.139000 0.458000 ;
        RECT 1.534000 0.530000 1.725000 0.585000 ;
        RECT 1.377000 0.650000 1.595000 0.705000 ;
        RECT 1.352000 0.287000 1.595000 0.342000 ;
        RECT 1.249000 0.520000 1.450000 0.575000 ;
        RECT 0.870000 0.265000 1.139000 0.320000 ;
        RECT 0.530000 0.995000 1.267000 1.050000 ;
        RECT 0.196000 0.812000 0.769000 0.867000 ;
        RECT 1.078000 0.404000 1.310000 0.458000 ;
        RECT 1.029000 0.779000 1.310000 0.833000 ;
        RECT 0.387000 0.236000 0.963000 0.290000 ;
    END
END AOI222X4

MACRO AOI222X2
    CLASS CORE ;
    FOREIGN AOI222X2 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 2.500000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.814000 0.556000 2.016000 0.627000 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 2.210000 0.439000 2.273000 0.545000 ;
        RECT 1.665000 0.439000 2.273000 0.494000 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.130000 0.558000 1.331000 0.627000 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.951000 0.439000 1.558000 0.494000 ;
        END
    END B1
    PIN C0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.319000 0.398000 0.517000 0.507000 ;
        END
    END C0
    PIN C1
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.628000 0.556000 0.725000 0.620000 ;
        RECT 0.093000 0.521000 0.156000 0.627000 ;
        RECT 0.093000 0.565000 0.299000 0.627000 ;
        RECT 0.093000 0.565000 0.725000 0.620000 ;
        END
    END C1
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 2.500000 1.280000 ;
        RECT 0.741000 0.911000 0.833000 1.280000 ;
        RECT 0.395000 0.911000 0.487000 1.280000 ;
        RECT 0.049000 0.911000 0.141000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 2.500000 0.080000 ;
        RECT 2.261000 -0.080000 2.353000 0.198000 ;
        RECT 1.567000 -0.080000 1.659000 0.198000 ;
        RECT 0.782000 -0.080000 0.874000 0.198000 ;
        RECT 0.049000 -0.080000 0.141000 0.275000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 2.263000 0.268000 2.399000 0.367000 ;
        RECT 1.905000 0.249000 2.024000 0.323000 ;
        RECT 1.190000 0.249000 1.318000 0.323000 ;
        RECT 2.336000 0.268000 2.399000 0.743000 ;
        RECT 2.201000 0.688000 2.263000 0.761000 ;
        RECT 1.797000 0.688000 2.399000 0.743000 ;
        RECT 0.395000 0.268000 2.399000 0.323000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.222000 0.688000 1.542000 0.743000 ;
        RECT 0.931000 0.910000 2.408000 0.964000 ;
    END
END AOI222X2

MACRO AOI222X1
    CLASS CORE ;
    FOREIGN AOI222X1 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.400000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.912000 0.444000 1.013000 0.627000 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.087000 0.433000 1.188000 0.587000 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.701000 0.433000 0.838000 0.535000 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.488000 0.506000 0.586000 0.627000 ;
        RECT 0.407000 0.573000 0.586000 0.627000 ;
        END
    END B1
    PIN C0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.037000 0.439000 0.122000 0.633000 ;
        END
    END C0
    PIN C1
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.232000 0.405000 0.380000 0.507000 ;
        END
    END C1
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 1.400000 1.280000 ;
        RECT 0.387000 0.917000 0.477000 1.280000 ;
        RECT 0.048000 0.941000 0.138000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 1.400000 0.080000 ;
        RECT 1.179000 -0.080000 1.269000 0.122000 ;
        RECT 0.418000 -0.080000 0.508000 0.122000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.282000 0.281000 1.343000 0.743000 ;
        RECT 1.083000 0.688000 1.343000 0.743000 ;
        RECT 0.048000 0.281000 1.343000 0.336000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.646000 0.685000 0.707000 0.817000 ;
        RECT 0.217000 0.762000 0.707000 0.817000 ;
        RECT 0.646000 0.685000 0.834000 0.739000 ;
        RECT 0.574000 0.910000 1.343000 0.964000 ;
    END
END AOI222X1

MACRO AOI221X4
    CLASS CORE ;
    FOREIGN AOI221X4 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 2.000000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.423000 0.433000 0.534000 0.585000 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.668000 0.502000 0.731000 0.627000 ;
        RECT 0.668000 0.567000 0.850000 0.627000 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.241000 0.598000 0.336000 0.761000 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.039000 0.462000 0.143000 0.632000 ;
        END
    END B1
    PIN C0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.862000 0.373000 1.032000 0.494000 ;
        END
    END C0
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 2.000000 1.280000 ;
        RECT 1.840000 0.765000 1.934000 1.280000 ;
        RECT 0.358000 1.078000 0.452000 1.280000 ;
        RECT 1.444000 0.765000 1.537000 1.280000 ;
        RECT 0.050000 1.078000 0.143000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 2.000000 0.080000 ;
        RECT 1.427000 -0.080000 1.521000 0.198000 ;
        RECT 0.766000 -0.080000 0.860000 0.122000 ;
        RECT 0.050000 -0.080000 0.143000 0.291000 ;
        RECT 1.843000 -0.080000 1.906000 0.361000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.675000 0.300000 1.780000 0.633000 ;
        RECT 1.642000 0.660000 1.738000 0.964000 ;
        RECT 1.675000 0.300000 1.738000 0.964000 ;
        RECT 1.625000 0.300000 1.780000 0.355000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 1.084000 0.723000 1.179000 0.810000 ;
        RECT 1.245000 0.895000 1.339000 0.976000 ;
        RECT 1.333000 0.345000 1.397000 0.644000 ;
        RECT 1.275000 0.589000 1.339000 0.976000 ;
        RECT 1.242000 0.274000 1.306000 0.400000 ;
        RECT 1.116000 0.236000 1.179000 0.810000 ;
        RECT 0.602000 0.236000 0.665000 0.306000 ;
        RECT 1.333000 0.508000 1.573000 0.563000 ;
        RECT 1.275000 0.589000 1.397000 0.644000 ;
        RECT 1.242000 0.345000 1.397000 0.400000 ;
        RECT 1.116000 0.468000 1.270000 0.523000 ;
        RECT 0.402000 0.251000 0.665000 0.306000 ;
        RECT 0.204000 0.832000 0.799000 0.887000 ;
        RECT 0.602000 0.236000 1.179000 0.290000 ;
        RECT 1.333000 0.345000 1.339000 0.976000 ;
    END
END AOI221X4

MACRO AOI221X2
    CLASS CORE ;
    FOREIGN AOI221X2 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 2.100000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.087000 0.396000 1.233000 0.500000 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.932000 0.573000 0.993000 0.650000 ;
        RECT 0.917000 0.595000 1.572000 0.650000 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.212000 0.306000 0.313000 0.430000 ;
        RECT 0.212000 0.375000 0.414000 0.430000 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.562000 0.433000 0.663000 0.558000 ;
        RECT 0.562000 0.493000 0.711000 0.558000 ;
        RECT 0.077000 0.504000 0.711000 0.558000 ;
        END
    END B1
    PIN C0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.678000 0.439000 1.739000 0.543000 ;
        RECT 1.457000 0.439000 1.739000 0.494000 ;
        END
    END C0
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 2.100000 1.280000 ;
        RECT 0.727000 0.903000 0.817000 1.280000 ;
        RECT 0.387000 0.903000 0.477000 1.280000 ;
        RECT 0.048000 0.903000 0.138000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 2.100000 0.080000 ;
        RECT 1.546000 -0.080000 1.636000 0.198000 ;
        RECT 0.780000 -0.080000 0.870000 0.122000 ;
        RECT 0.048000 -0.080000 0.138000 0.198000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.761000 0.755000 1.868000 0.836000 ;
        RECT 1.330000 0.300000 1.457000 0.367000 ;
        RECT 1.807000 0.312000 1.868000 0.836000 ;
        RECT 1.330000 0.225000 1.391000 0.367000 ;
        RECT 1.330000 0.312000 1.868000 0.367000 ;
        RECT 0.387000 0.225000 1.391000 0.280000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.883000 0.707000 0.944000 0.823000 ;
        RECT 0.912000 0.962000 2.020000 1.017000 ;
        RECT 0.883000 0.768000 1.511000 0.823000 ;
        RECT 0.217000 0.707000 0.944000 0.762000 ;
    END
END AOI221X2

MACRO AOI221X1
    CLASS CORE ;
    FOREIGN AOI221X1 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.300000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.432000 0.306000 0.560000 0.431000 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.803000 0.379000 0.868000 0.494000 ;
        RECT 0.667000 0.379000 0.868000 0.433000 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.225000 0.520000 0.380000 0.633000 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.049000 0.306000 0.146000 0.461000 ;
        END
    END B1
    PIN C0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.979000 0.393000 1.044000 0.627000 ;
        RECT 0.979000 0.573000 1.054000 0.627000 ;
        END
    END C0
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 1.300000 1.280000 ;
        RECT 0.411000 0.916000 0.506000 1.280000 ;
        RECT 0.051000 0.916000 0.146000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 1.300000 0.080000 ;
        RECT 0.782000 -0.080000 0.878000 0.122000 ;
        RECT 0.051000 -0.080000 0.146000 0.229000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.165000 0.627000 1.240000 0.754000 ;
        RECT 0.632000 0.227000 0.703000 0.312000 ;
        RECT 1.175000 0.257000 1.240000 0.761000 ;
        RECT 0.632000 0.189000 0.696000 0.312000 ;
        RECT 0.632000 0.257000 1.240000 0.312000 ;
        RECT 0.411000 0.189000 0.696000 0.244000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.609000 0.862000 1.065000 0.917000 ;
        RECT 0.231000 0.689000 0.885000 0.744000 ;
    END
END AOI221X1

MACRO AOI21XL
    CLASS CORE ;
    FOREIGN AOI21XL 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 0.700000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.212000 0.567000 0.379000 0.662000 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.045000 0.417000 0.138000 0.562000 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.362000 0.411000 0.513000 0.500000 ;
        END
    END B0
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 0.700000 1.280000 ;
        RECT 0.223000 1.078000 0.313000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 0.700000 0.080000 ;
        RECT 0.536000 -0.080000 0.626000 0.122000 ;
        RECT 0.048000 -0.080000 0.138000 0.331000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.582000 0.295000 0.643000 0.627000 ;
        RECT 0.573000 0.573000 0.634000 0.830000 ;
        RECT 0.387000 0.295000 0.643000 0.350000 ;
        RECT 0.573000 0.573000 0.643000 0.627000 ;
        RECT 0.582000 0.295000 0.634000 0.830000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.374000 0.952000 0.435000 1.050000 ;
        RECT 0.062000 0.749000 0.123000 1.007000 ;
        RECT 0.374000 0.995000 0.498000 1.050000 ;
        RECT 0.062000 0.952000 0.435000 1.007000 ;
    END
END AOI21XL

MACRO AOI21X4
    CLASS CORE ;
    FOREIGN AOI21X4 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.800000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.115000 0.469000 0.207000 0.574000 ;
        RECT 0.745000 0.530000 0.807000 0.627000 ;
        RECT 0.145000 0.469000 0.207000 0.625000 ;
        RECT 0.145000 0.567000 0.218000 0.625000 ;
        RECT 0.145000 0.570000 0.807000 0.625000 ;
        RECT 0.745000 0.573000 0.841000 0.627000 ;
        RECT 0.145000 0.573000 0.841000 0.625000 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.415000 0.392000 0.661000 0.494000 ;
        RECT 1.005000 0.452000 1.098000 0.533000 ;
        RECT 0.400000 0.426000 0.492000 0.507000 ;
        RECT 0.415000 0.392000 0.492000 0.507000 ;
        RECT 0.400000 0.426000 0.661000 0.494000 ;
        RECT 1.005000 0.392000 1.068000 0.533000 ;
        RECT 0.415000 0.392000 1.068000 0.446000 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.238000 0.496000 1.402000 0.635000 ;
        END
    END B0
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 1.800000 1.280000 ;
        RECT 0.922000 0.941000 1.015000 1.280000 ;
        RECT 0.573000 0.941000 0.665000 1.280000 ;
        RECT 0.224000 0.941000 0.316000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 1.800000 0.080000 ;
        RECT 1.458000 -0.080000 1.550000 0.122000 ;
        RECT 1.098000 -0.080000 1.190000 0.198000 ;
        RECT 0.400000 -0.080000 0.492000 0.198000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.208000 0.274000 1.319000 0.392000 ;
        RECT 1.478000 0.300000 1.582000 0.633000 ;
        RECT 1.620000 0.896000 1.713000 0.977000 ;
        RECT 1.271000 0.896000 1.364000 0.977000 ;
        RECT 1.605000 0.896000 1.713000 0.964000 ;
        RECT 1.605000 0.579000 1.668000 0.964000 ;
        RECT 1.208000 0.337000 1.582000 0.392000 ;
        RECT 0.049000 0.274000 1.319000 0.329000 ;
        RECT 1.478000 0.579000 1.668000 0.633000 ;
        RECT 1.271000 0.910000 1.713000 0.964000 ;
        RECT 1.620000 0.579000 1.668000 0.977000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.049000 0.698000 1.538000 0.752000 ;
    END
END AOI21X4

MACRO AOI21X1
    CLASS CORE ;
    FOREIGN AOI21X1 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 0.700000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.232000 0.306000 0.293000 0.623000 ;
        RECT 0.232000 0.568000 0.379000 0.623000 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.050000 0.492000 0.141000 0.615000 ;
        RECT 0.050000 0.433000 0.138000 0.615000 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.477000 0.439000 0.542000 0.627000 ;
        RECT 0.407000 0.439000 0.542000 0.494000 ;
        END
    END B0
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 0.700000 1.280000 ;
        RECT 0.217000 0.852000 0.308000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 0.700000 0.080000 ;
        RECT 0.536000 -0.080000 0.626000 0.122000 ;
        RECT 0.048000 -0.080000 0.138000 0.334000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.582000 0.706000 0.664000 0.940000 ;
        RECT 0.387000 0.295000 0.477000 0.376000 ;
        RECT 0.557000 0.860000 0.664000 0.940000 ;
        RECT 0.603000 0.321000 0.664000 0.940000 ;
        RECT 0.387000 0.321000 0.664000 0.376000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.048000 0.696000 0.477000 0.751000 ;
    END
END AOI21X1

MACRO AND4XL
    CLASS CORE ;
    FOREIGN AND4XL 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.100000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.039000 0.606000 0.144000 0.767000 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.222000 0.508000 0.328000 0.688000 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.406000 0.508000 0.511000 0.688000 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.706000 0.573000 0.863000 0.688000 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.258000 1.078000 0.861000 1.280000 ;
        RECT 0.000000 1.120000 1.100000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 1.100000 0.080000 ;
        RECT 0.739000 -0.080000 0.833000 0.122000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.950000 0.760000 1.061000 0.900000 ;
        RECT 0.965000 0.242000 1.029000 0.900000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.533000 0.751000 0.628000 0.887000 ;
        RECT 0.575000 0.367000 0.896000 0.455000 ;
        RECT 0.050000 0.232000 0.144000 0.313000 ;
        RECT 0.533000 0.751000 0.639000 0.824000 ;
        RECT 0.575000 0.232000 0.639000 0.824000 ;
        RECT 0.144000 0.832000 0.628000 0.887000 ;
        RECT 0.050000 0.232000 0.639000 0.287000 ;
        RECT 0.575000 0.232000 0.628000 0.887000 ;
    END
END AND4XL

MACRO AND4X4
    CLASS CORE ;
    FOREIGN AND4X4 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 2.000000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.579000 0.625000 0.689000 0.773000 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.766000 0.489000 0.871000 0.629000 ;
        RECT 0.460000 0.489000 0.871000 0.544000 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.220000 0.493000 0.344000 0.636000 ;
        RECT 0.220000 0.539000 0.364000 0.636000 ;
        RECT 0.988000 0.379000 1.051000 0.721000 ;
        RECT 0.281000 0.379000 0.344000 0.636000 ;
        RECT 0.948000 0.379000 1.051000 0.439000 ;
        RECT 0.281000 0.379000 1.051000 0.433000 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.039000 0.640000 0.146000 0.767000 ;
        RECT 1.213000 0.567000 1.328000 0.650000 ;
        RECT 1.264000 0.439000 1.328000 0.650000 ;
        RECT 1.114000 0.595000 1.178000 0.888000 ;
        RECT 0.081000 0.640000 0.145000 0.888000 ;
        RECT 1.264000 0.439000 1.364000 0.494000 ;
        RECT 1.114000 0.595000 1.328000 0.650000 ;
        RECT 0.081000 0.833000 1.178000 0.888000 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 2.000000 1.280000 ;
        RECT 1.643000 1.078000 1.751000 1.280000 ;
        RECT 0.251000 1.078000 0.358000 1.280000 ;
        RECT 1.131000 1.078000 1.225000 1.280000 ;
        RECT 0.689000 1.078000 0.782000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 2.000000 0.080000 ;
        RECT 1.372000 -0.080000 1.466000 0.250000 ;
        RECT 1.769000 -0.080000 1.862000 0.211000 ;
        RECT 0.050000 -0.080000 0.143000 0.334000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.675000 0.567000 1.780000 0.900000 ;
        RECT 1.438000 0.815000 1.532000 1.039000 ;
        RECT 1.438000 0.815000 1.780000 0.900000 ;
        RECT 1.676000 0.356000 1.759000 0.900000 ;
        RECT 1.675000 0.356000 1.759000 0.439000 ;
        RECT 1.570000 0.331000 1.696000 0.412000 ;
        RECT 1.570000 0.356000 1.759000 0.412000 ;
        RECT 1.676000 0.331000 1.696000 0.900000 ;
        RECT 1.675000 0.331000 1.676000 0.439000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.905000 0.944000 0.999000 1.039000 ;
        RECT 0.479000 0.944000 0.573000 1.039000 ;
        RECT 1.444000 0.507000 1.574000 0.588000 ;
        RECT 0.711000 0.240000 0.804000 0.321000 ;
        RECT 1.242000 0.706000 1.306000 0.999000 ;
        RECT 1.444000 0.329000 1.507000 0.761000 ;
        RECT 1.164000 0.254000 1.227000 0.383000 ;
        RECT 1.242000 0.706000 1.507000 0.761000 ;
        RECT 0.479000 0.944000 1.306000 0.999000 ;
        RECT 1.164000 0.329000 1.507000 0.383000 ;
        RECT 0.905000 0.254000 1.227000 0.308000 ;
        RECT 0.804000 0.254000 1.164000 0.308000 ;
        RECT 0.711000 0.254000 0.999000 0.308000 ;
    END
END AND4X4

MACRO AND4X2
    CLASS CORE ;
    FOREIGN AND4X2 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.100000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.039000 0.398000 0.157000 0.556000 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.222000 0.537000 0.358000 0.645000 ;
        RECT 0.279000 0.537000 0.358000 0.646000 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.478000 0.581000 0.542000 0.761000 ;
        RECT 0.426000 0.706000 0.542000 0.761000 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.610000 0.439000 0.694000 0.606000 ;
        RECT 0.610000 0.524000 0.733000 0.606000 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 1.100000 1.280000 ;
        RECT 0.724000 1.064000 0.838000 1.280000 ;
        RECT 0.049000 1.078000 0.158000 1.280000 ;
        RECT 0.419000 1.078000 0.514000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 1.100000 0.080000 ;
        RECT 0.721000 -0.080000 0.815000 0.122000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.967000 0.648000 1.049000 0.767000 ;
        RECT 0.967000 0.700000 1.061000 0.767000 ;
        RECT 0.985000 0.358000 1.049000 0.767000 ;
        RECT 0.967000 0.648000 1.031000 0.964000 ;
        RECT 0.967000 0.199000 1.031000 0.413000 ;
        RECT 0.967000 0.358000 1.049000 0.413000 ;
        RECT 0.985000 0.199000 1.031000 0.964000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.061000 0.250000 0.156000 0.343000 ;
        RECT 0.825000 0.473000 0.919000 0.556000 ;
        RECT 0.076000 0.211000 0.156000 0.343000 ;
        RECT 0.825000 0.211000 0.889000 0.889000 ;
        RECT 0.208000 0.835000 0.889000 0.889000 ;
        RECT 0.076000 0.211000 0.889000 0.265000 ;
    END
END AND4X2

MACRO AND4X1
    CLASS CORE ;
    FOREIGN AND4X1 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.100000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.039000 0.615000 0.147000 0.776000 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.175000 0.399000 0.328000 0.545000 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.392000 0.567000 0.511000 0.696000 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.703000 0.573000 0.857000 0.696000 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.258000 1.078000 0.861000 1.280000 ;
        RECT 0.000000 1.120000 1.100000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 1.100000 0.080000 ;
        RECT 0.739000 -0.080000 0.833000 0.122000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.956000 0.761000 1.061000 0.905000 ;
        RECT 0.950000 0.800000 1.061000 0.905000 ;
        RECT 0.950000 0.244000 1.044000 0.325000 ;
        RECT 0.981000 0.244000 1.044000 0.905000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.533000 0.751000 0.628000 0.887000 ;
        RECT 0.814000 0.401000 0.908000 0.482000 ;
        RECT 0.050000 0.223000 0.144000 0.304000 ;
        RECT 0.533000 0.751000 0.639000 0.824000 ;
        RECT 0.814000 0.223000 0.878000 0.482000 ;
        RECT 0.575000 0.414000 0.639000 0.824000 ;
        RECT 0.575000 0.414000 0.908000 0.469000 ;
        RECT 0.144000 0.832000 0.628000 0.887000 ;
        RECT 0.050000 0.223000 0.878000 0.277000 ;
        RECT 0.575000 0.414000 0.628000 0.887000 ;
    END
END AND4X1

MACRO AND3XL
    CLASS CORE ;
    FOREIGN AND3XL 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 0.900000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.038000 0.426000 0.158000 0.548000 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.172000 0.677000 0.310000 0.786000 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.397000 0.408000 0.539000 0.511000 ;
        END
    END C
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 0.900000 1.280000 ;
        RECT 0.273000 1.078000 0.365000 1.280000 ;
        RECT 0.610000 0.639000 0.734000 0.729000 ;
        RECT 0.275000 1.065000 0.364000 1.280000 ;
        RECT 0.610000 0.639000 0.672000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 0.900000 0.080000 ;
        RECT 0.545000 -0.080000 0.638000 0.122000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.747000 0.832000 0.862000 1.010000 ;
        RECT 0.758000 0.274000 0.859000 0.355000 ;
        RECT 0.796000 0.274000 0.859000 1.010000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.055000 0.940000 0.147000 1.037000 ;
        RECT 0.633000 0.417000 0.734000 0.500000 ;
        RECT 0.049000 0.255000 0.142000 0.336000 ;
        RECT 0.400000 0.567000 0.477000 0.744000 ;
        RECT 0.225000 0.268000 0.288000 0.621000 ;
        RECT 0.633000 0.268000 0.695000 0.500000 ;
        RECT 0.415000 0.567000 0.477000 0.995000 ;
        RECT 0.147000 0.268000 0.695000 0.323000 ;
        RECT 0.055000 0.940000 0.477000 0.995000 ;
        RECT 0.049000 0.268000 0.477000 0.323000 ;
        RECT 0.225000 0.567000 0.477000 0.621000 ;
    END
END AND3XL

MACRO AND2XL
    CLASS CORE ;
    FOREIGN AND2XL 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 0.700000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.040000 0.433000 0.150000 0.551000 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.219000 0.564000 0.320000 0.702000 ;
        END
    END B
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.122000 1.078000 0.371000 1.280000 ;
        RECT 0.000000 1.120000 0.700000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 0.700000 0.080000 ;
        RECT 0.384000 -0.080000 0.475000 0.122000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.563000 0.567000 0.663000 0.633000 ;
        RECT 0.563000 0.344000 0.624000 0.845000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.048000 0.182000 0.138000 0.263000 ;
        RECT 0.122000 0.760000 0.212000 0.840000 ;
        RECT 0.440000 0.195000 0.501000 0.827000 ;
        RECT 0.212000 0.195000 0.501000 0.250000 ;
        RECT 0.138000 0.195000 0.440000 0.250000 ;
        RECT 0.048000 0.195000 0.212000 0.250000 ;
        RECT 0.122000 0.773000 0.501000 0.827000 ;
    END
END AND2XL

MACRO AND2X4
    CLASS CORE ;
    FOREIGN AND2X4 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 0.900000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.038000 0.482000 0.142000 0.660000 ;
        RECT 0.038000 0.482000 0.145000 0.574000 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.218000 0.627000 0.322000 0.786000 ;
        RECT 0.312000 0.471000 0.375000 0.562000 ;
        RECT 0.259000 0.507000 0.322000 0.786000 ;
        RECT 0.259000 0.507000 0.375000 0.562000 ;
        RECT 0.312000 0.471000 0.322000 0.786000 ;
        END
    END B
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 0.900000 1.280000 ;
        RECT 0.046000 1.078000 0.146000 1.280000 ;
        RECT 0.755000 0.914000 0.848000 1.280000 ;
        RECT 0.394000 1.078000 0.487000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 0.900000 0.080000 ;
        RECT 0.755000 -0.080000 0.848000 0.243000 ;
        RECT 0.387000 -0.080000 0.480000 0.122000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.592000 0.326000 0.784000 0.433000 ;
        RECT 0.758000 0.433000 0.862000 0.767000 ;
        RECT 0.758000 0.331000 0.860000 0.798000 ;
        RECT 0.592000 0.331000 0.860000 0.433000 ;
        RECT 0.580000 0.717000 0.860000 0.798000 ;
        RECT 0.580000 0.717000 0.862000 0.767000 ;
        RECT 0.758000 0.326000 0.784000 0.798000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.440000 0.498000 0.663000 0.579000 ;
        RECT 0.049000 0.343000 0.142000 0.424000 ;
        RECT 0.440000 0.354000 0.503000 0.671000 ;
        RECT 0.386000 0.617000 0.449000 0.910000 ;
        RECT 0.202000 0.855000 0.449000 0.910000 ;
        RECT 0.386000 0.617000 0.503000 0.671000 ;
        RECT 0.202000 0.354000 0.503000 0.408000 ;
        RECT 0.142000 0.354000 0.440000 0.408000 ;
        RECT 0.049000 0.354000 0.386000 0.408000 ;
        RECT 0.440000 0.354000 0.449000 0.910000 ;
    END
END AND2X4

MACRO AND2X2
    CLASS CORE ;
    FOREIGN AND2X2 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 0.700000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.037000 0.504000 0.138000 0.633000 ;
        RECT 0.037000 0.504000 0.202000 0.585000 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.212000 0.833000 0.361000 0.935000 ;
        END
    END B
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 0.700000 1.280000 ;
        RECT 0.048000 1.078000 0.151000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 0.700000 0.080000 ;
        RECT 0.350000 -0.080000 0.440000 0.122000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.552000 0.227000 0.654000 0.390000 ;
        RECT 0.552000 0.688000 0.642000 1.002000 ;
        RECT 0.552000 0.195000 0.642000 0.390000 ;
        RECT 0.552000 0.688000 0.654000 0.767000 ;
        RECT 0.582000 0.227000 0.654000 0.439000 ;
        RECT 0.593000 0.227000 0.654000 0.767000 ;
        RECT 0.582000 0.195000 0.642000 0.439000 ;
        RECT 0.593000 0.195000 0.642000 1.002000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.216000 0.654000 0.325000 0.737000 ;
        RECT 0.264000 0.512000 0.521000 0.594000 ;
        RECT 0.048000 0.321000 0.138000 0.402000 ;
        RECT 0.264000 0.348000 0.325000 0.737000 ;
        RECT 0.048000 0.348000 0.325000 0.402000 ;
    END
END AND2X2

MACRO AND2X1
    CLASS CORE ;
    FOREIGN AND2X1 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 0.700000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.040000 0.433000 0.150000 0.551000 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.212000 0.551000 0.322000 0.689000 ;
        END
    END B
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 0.700000 1.280000 ;
        RECT 0.347000 1.078000 0.465000 1.280000 ;
        RECT 0.119000 1.078000 0.209000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 0.700000 0.080000 ;
        RECT 0.384000 -0.080000 0.475000 0.122000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.549000 0.732000 0.639000 0.927000 ;
        RECT 0.549000 0.320000 0.639000 0.401000 ;
        RECT 0.562000 0.320000 0.639000 0.439000 ;
        RECT 0.563000 0.567000 0.663000 0.633000 ;
        RECT 0.563000 0.320000 0.624000 0.927000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.048000 0.182000 0.138000 0.263000 ;
        RECT 0.119000 0.760000 0.209000 0.840000 ;
        RECT 0.423000 0.461000 0.500000 0.561000 ;
        RECT 0.426000 0.195000 0.487000 0.827000 ;
        RECT 0.209000 0.195000 0.487000 0.250000 ;
        RECT 0.138000 0.195000 0.426000 0.250000 ;
        RECT 0.048000 0.195000 0.423000 0.250000 ;
        RECT 0.119000 0.773000 0.487000 0.827000 ;
    END
END AND2X1

MACRO BUFX6
    CLASS CORE ;
    FOREIGN BUFX6 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.300000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.160000 0.474000 0.391000 0.555000 ;
        RECT 0.246000 0.439000 0.311000 0.555000 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 1.300000 1.280000 ;
        RECT 0.422000 1.078000 0.518000 1.280000 ;
        RECT 1.154000 0.877000 1.249000 1.280000 ;
        RECT 0.794000 0.877000 0.889000 1.280000 ;
        RECT 0.051000 0.844000 0.146000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 1.300000 0.080000 ;
        RECT 0.816000 -0.080000 0.912000 0.215000 ;
        RECT 0.456000 -0.080000 0.552000 0.215000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.803000 0.433000 1.240000 0.767000 ;
        RECT 0.803000 0.321000 1.126000 0.767000 ;
        RECT 0.782000 0.625000 1.240000 0.757000 ;
        RECT 0.782000 0.321000 1.126000 0.440000 ;
        RECT 0.636000 0.321000 1.126000 0.402000 ;
        RECT 0.613000 0.676000 1.240000 0.757000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.484000 0.519000 0.718000 0.600000 ;
        RECT 0.253000 0.274000 0.349000 0.355000 ;
        RECT 0.231000 0.657000 0.326000 0.738000 ;
        RECT 0.484000 0.300000 0.549000 0.712000 ;
        RECT 0.253000 0.300000 0.549000 0.355000 ;
        RECT 0.231000 0.657000 0.549000 0.712000 ;
    END
END BUFX6

END LIBRARY
